%PDF-1.7

4 0 obj
(Identity)
endobj
5 0 obj
(Adobe)
endobj
8 0 obj
<<
/Filter /FlateDecode
/Length 67006
/Length1 325580
/Type /Stream
>>
stream
x��`\U���y͙�#3��L���$i�I2y?ڴ�&Mߥ����M��I�)�R�H}`1����"rQQd����B�V.
U^�PA@D\E�B�����Ʉ��^�����Yg�}��g���^k��� ?	�f-�7玚�V��(88gV��;7�Ħ��9K/��i�^���Q=gي�������\v�������k�<
���{��e��_w�x���O��g�SWt,_ ?����C��/�-��?�~�ȧ���@��8��n�t�[f>���+�ڋ����y�z��K7V_��}`�3����w��� +�@ݲy�ځW?68�����͘�1��
���ś�߱��g@�H~�^���>���n[��g��]5���+������|s=��?��G�߰c���F�@��r<�u���7���N���G��]�#���~�^?tᆡ-G~k�X_���&��;��k�m��
?9�O������Né�����h��T2�������e��YIYp�Bs��a�X���$|��'+D�3�:�A��"�c�%�^�>&�SA�*�(K� =���_����-�D���;�R�u����!�H�H��0}S�S�*	{��=�	.��%Dg�e�\X��󸝏�Z��pۍ�
���6�N�1���#=�~�H����p�?z�R7��h�H[����a���tzB����{n�u����� \-�i��&5�4�O�;�j�\���K_���i���FY��x���=� �ۃ�*��P�ߧ���Ц���*���������������������������������������� �;l��5�W���������������0�
������� &�j��dP�� 8-�ـʀ�C�.>����6[�
PY�E`���؀����������gΰ����?� ppLh��Il��������V�"��==
vF�L�'��������A�>�^�E�?�\F���~� �~E�� ���� i>"-`�"H�EA�_�"�EP�4%H��i	LI��P�t
�eP��;�CiT"�C�J�N�	U�VC��"��:��P����C���FhF�-H�m�i�7�ڐN��H�1�3�N�v�3 ��+����_ 	�Hg2���v�l��`�.Fg�\�s`>ҹ� ��0�_����F�YH�b�g��H�R�K`ҳay�5X��2�F��A���n�M�
��J�=�*}za5ҕЇt��t5�?C�Az.�C���~X�t-���]��&�`ҍH_�M��fD��ѭp>�����a���a;��B���"�CH_��酰�Ep	�p)ҋ��K���K�r���
���G�^��E��D�>��
�ҏ�Ǒ^	�H��0�Q�
����H?�B�	�/�U0���pҽ�^�F�)�L��0��5p�k�sH?ק���0�Y�����H?������×����"|��Ho�����5�_���~nA�UFo�C�5�f�wp3�_�[���B�o�m��@�|���V��������������w�N��C*�[��߇}H�H ���h
!�w��= G���H��!�;�k��!=�"=��QAz7�{�)8���'H���{�>�#�H��G�c�ҟ�ϑ���L?�1�����p?<��g��F� <��Ax�	x�/�q���'ҿ��}�D�<��Q�5���7���W�4����O }��g�>�!�5����ӏ�o��H��? }^D�;x	��2��}^A�{�S�ax���p��*җ�>/��H������?1�gx�Ix3�Kx�/�5�;���-����_�m��SH�`�o0��MK���C�[����m" }��HO	�(Q��1�&&��zܛ�f3�"Hي_�3��)�Y�
(
=��dY�)@TL�(�����ĢO�����������C�3
�I��8]0�d�b��'�"��Y�����Y2�
��LA��$ITX�E���MǙ �(p'���tA�ɂ�j}o�E����,��8�Ȋ��,�g�%g����������q�MIs'���t��Y8&6�$ib0D6e��YT^�`V�ޙLTl�,(&�D3�z���b��ə��&���������L ��ppp�S0�d�n���8���g��8����	��gA�4�"+Ҥ�YD���������������N*��88&���Y&Cd5��8��0r3���,*�T��*�I��S���X�-}�I �*��������8��,����1Yp:� ��,�{�,�8����,�,�RAUM���Y�,�b�q�g��g��8]��d��r�7�b�@Ϸ�a�lV�wsV����dV�l�@�f�VL�Y����LBL�&�����������2ΰ��<���q���,���M�,���/�b3����Y�,΢g��lV��	qU1�vg����������W��,����1Y�x<�(X2x�8�Æ��j����Y0[T�,	̒�baq��N#0��ؓ�Y88888888��a?���T��ppLrrrh�e¢��8���e,�v���j��ݳ��j�Z�j�q���*V���Y888888888��8�?'ppL�^�{�,�5=�bpd�Y�`�� �ɛ�V��R,���`Lf�����Y�)Ǉg�O,�8����pL|>�L�]���>��r����&�Yl�l6g�`��0����q�<�����O�����\g��q�j�@������s;��9lv����l6����,V�CC0��d��hfr{�8Ǚ�3�,y����t������8�ٞ�gq �#�q��sس�,v�٭v��4Βcgq�nu�8ǿ�3�,����q����B^^��ď{�q�%�vp���{v�ۭv;���d/������+]&g�'7agx�����BppLB���LXtbqf��_\l����v� �ɛN��N�v���+-6�����Y� Ǉg�O,�8��88&`6O\tbue��Y� ^���栽�ܐ���N�����S����-.G.8ؿI�	888888888>�8�~b�Orp�.��d!���2qщ͝���%����-�x=9�Y�����q��c�)�)�9�W��L�����,gΰ��<���q� ��B4}O����@_��e�X4r�g�d�,*��|���z\p�� 888888888>���>��q���,������&.:qx3��/�l��� �;��.�ҳ���u{s��S���}h�n���7	�q�3g��g��8]( ��BEE���|u�3��/��<�l$�����\�?�~�,1����������LBX����������Ï3lJ�Orp�.D��c�P]]��E'�@�G?� �~6F{Wa2�� /��A h�uJ͡����hfr&!������������G�(������ ����:p�&.:�	e��_
����S���|�K_��`�??��VX+��zr����1��^�8Ǚ�B8��]sp�.L��BSS����
2��6Pb��b�wE�tVX�)���@a>� d�*, �����h�0	�Ǉg��>��q�P���S������H�/���2US��G�0Y��D�0��!�C��6���̉�i�a`�?������8]���Bgg'�|�|�d��S�bZ��m���(�˰��X%+	�Ġ��	QgKI1@^anI����I'ppppppppp|�Qg�d ��BppL,X ~��/_�3��/U �ƺ��uP��JLVj9�0�<V>�+�P�n�(E%-P��o��?ΰ)i>��q�088&˖-�`��y���_��hI�g��P�5���r��������s�<gv5�����Pe�3	�~��>��q������ի�� J��bu��f�ƺ�9ӡZ�0٨��AM}E}����ڷ�� Z����Pi,z9��Ǉ�pF��s��c�000 ���E'�����x����N�w3Z�2,})V344W77Bs����[� ���-u�i�X�rz��?��/ppp�,�I7���܏�j�`ʁ���L肳`	,�X`l�K�R���[Hm�\��;J:��O���P���Rv�Z�����>������������r�g��_ ��]�}h����u��M7�[sn��U+{{V,_���%���9�{��mӦ��4756����$��*��eSJK�cE�H�� ?��s}����t�mV�Y5)�$
*I*��g_�E���*�88�8%���M�g�E�wݔ���wf��J�75;�9��f�����>��,�'�7ul�umI:���Y1W$5���^V�>��3ֹ�RU	�,VLZ1���#�g�fwM�'�j��Ly�)���n[S�k�1��%ᙜ�3��#�f���H�h)�R:S&��ȖTrm
���������m�����sk���@,�ڼ��n��#)	g$�9��͑�eG��~��Yx���cvng���H(��}W�O��+�\�BH�������{#�[���>����7+<�������*y��J�t�o��ܺ�ֳkkd����ײ:�K�6cì����u���J�L%��,_��^Y7�W��/�3;�?�7�1{�ҞNZ���Y!��39�zft'#��Td}$K{bxi%Z`x}�h/����ߕ�K\���� E�c'�<1g������49;6�xxv,2{�x����u��+6�o��ᡮ~|���p��5���k{S���d*�J��=���8\b�
���r���;�2,�F�Q+zzCȧ�^�imO	��Xg�ц�{:�d4J���IX��=g�h�X��Dۣ��1��V�3{�3���c���L��Rji�������<5Er�����TNg�z��i�Ǟޖ��1]�Fx(�r�Sr�H��7�r����,���=���h9��R9@Q���<�w%*�`��p*�إ�A��Y����^K�Otؕ��f4v�<����й�'���b�K����*�^��#W��/I�^�������{�D�����W��z�D�$�\���Lz���v���ʮI�ag%����&��T#���Â���T���Hڙ�q��y���G��L�Z�3.z�(�=vR�>��IZ䤚4'm�]�#4k?��k�؈���a�KY�a�g�9Ү؃W$��_�b�b+V����(>��Bo	�0�`YJ*����,�rN�����S$�Z��uOu�.�bf,���������������;����(=E*�^��P~o,�І�2}p �v���.7�v!>�&��ǥֿ�Ӱ�)��R�Ǫ��	b��R��ë�WƢ�h��>X�:�{Y	X�YMbTUP#�&*���r�5���q|�uq,�gVl���������^�: S���I��6S-7�70[��ҕ���hx��.��r��r����'K�1oO&k>�=XA���q��ی��'���Kzv�n��.�jZ��D΀���5Vl)KlCG����4�]�Wh�)ց
�p�Z���Z����BE�ąZ��N��l��썢�\��ws�7��u>^7�n��='�g�ZZ�o�^Sɼ��)5S ^2/e��z	x�lv����(kkc,������M���C{��"W
�Ʀ��R�L��>(�;��1�N)IYJ�ҝ�hXN�a��L6����Z��ddYOT����l�Q7���O}-��j����X �Ѵ��?So�Vyv�W� ��JY�F�Y��o@��y�.���J/�wZ�هail�sZiV�	O���H�6��bN�Ÿ�RY-㸖k�onC��J8��6��,��~�?�_���yWFj�p�ݹv�=<�����_�=�g�B��T�#��1y���'�g{�����x�t[;���D#���uɨ���H�E�I`���GD?Қq8�i�����l����Uk.�s����� ʤq	m���T�<Ne7ϡ[?6O�C�ࣼ��g}�g������=<�z�ku��OJ]�P$��b���I�Y�����J�F��~���Ƶ�dl-5K��Y�~��S�j\B)���n��D�z{5��:Jz����p-�p��b,�;�<�ÿ�xl�lE�������X]�ZZ�+��xf3^"�P魣d�pK��G/��=������C�!����G#EmQ�5��!�ѣ^,H��\B/Ԅ������>S�x���.VY�l��Zb\�zMl�Ѣ�Oҗ'K٘�i(�����M�T���h�뾥v�<zk�h0�6��5<w�Y�J��K����g��U!dlվ�0�C�@S�B���:�Dh'���ģ$�v���)y�l��5&��S�����xg�%���u����w�)�Dڎ�ܮ�MJ��e����`b�~OK����AO�b�gh�;DV�k�	���A���|>���r�;z�-4cH���=ѷߧ%������ܥFb��D��p�����f;K�5��7鉲
=Q�Jn���K���3�]O��=�ê����N�k��ձ��w��Z�5���%��-##�����M  �.�z�4E���ޟ�m���z�A�ݔ��1aq����y,1}���$�ֺ�K/�_~�&9FZ�[����b^x��L#u��0iƽ���n�7��i�cB�H=80��^�ג���p�(iAjI�%8����z�����)��Sd�)���G�-���%=JF��?�~��`xϯȯp~�=A~��������sb���E���nZ��d2����ɵ?�?�����{�߲?������}�p������m:�~��AW��&�Φ����. �ngŘo�³�=����yȃ��[��^`�4}�$7�mC�l�ecj�t�{7��$+�m�_y���:2�r�_�V�s�uK֍��k��
�U�U׭��#޺�f���ܪ��p��$���+�9�ߕ�V&�����2�+|s�3��qt�x��_.Cs¡`[8�����̰��q�wfg(�I�/A��6r%���K~I^#ibqqB�a\	w½�Kx�`����N�)
�~)���(�쭲�*
�Z�%Kdr�Gm�g�r�u�˭�/H,��ӟ.�H}�:��=���.@��g�٢�`��8��wю�ؕR�6�E�o�E��A�Y�H9i��ERޮ�)olV��x6�=�#N��NA���ά���ggw�[X�b�
��ފ�{����^���/�������=��{~�=�4|�Hy��#u�øil&%��ׅ�p��>=<�=�l/w�/��-�[{c]��~ \��nlXnh,?��l���������B�̋�<-lQ���T/�q�Wb��ܱc�A�K��aȎ��v�1>�ںk3d8��>�B�+�.?,���G��C���sc���zů����Kp;����@�1�1���0L2� ����k-7���=Ha�L]A6��p˽�?�p~�߆�%��u�O/�j�G�	���g����ݗu�հZ��?����J�A�S�6A�b@��nD|D�6,�#�8��>7���/�@���|Q��߆��>�÷�m���Y�*���[�a�-�eB�a������q���)'?��
�@�r�~����?�\�ȭ/'�ᘐ�$#�Cy{[����b�"6���m���+��עd�Ϡ|Pl�_������x��p�x�X���tXG.'*��
����<��C�ܞ'?A���1،�vL��)��gXg�v;�K:$�
>��v)p�	}4�&�ޥ�-q�����D�Qw	�W��G�w�0����/�{j�xO�+(
�T��T	&�)bM��������V�h��	�P�&��x}�xMm/c�p<���͸)��	�t�B���1�I��&�"��A�
�(�$B�B�>��ښ�ru|��C��>"A�'1"<9z��,���wL=�����IV�5�B���r}d���̷^斧���}]Q�|8�z2��i��R��="Z�w���{�$�4w;�.4.N?v�n�a���6K<~�je�g1G�v;K��S���J��^��$�Uѫ`��~Y{�!L�lV�a|��;�EQ�f�c��n�f��	�H���P\�J.� �Z�F/Ez8�<{4&F���Jb\q����'����d�IL�����6���1zdP� {��q�`�+�.O}��4556�N)-�)&E�ys����uM���}�E��� /��p��e�ss"�u/;O��ض�O�������ⱏ�:4���|��/>k�˟��e��-��ϣ��G&c��)�Y����&�܉���VA����U玫۪R�X#$"�A	B��&ƒVzJ�Q�����h"���'����Ӫs���$ݵ�QD�����<�T�C��rD<<�=�uOR�E��ث뚚��Q��hq���˟3��7�/^}Υo������S$�u(�ﲷ�����x�Mn��ʳ��b��+���6��C;���.�\Y���:���(Q�\�����Ru\fC�j�=q���/��[���ʊ���x,�f!���O$t��7�kǎ�����G����ju�x��jMM���ü��\���_T�NmY�Z~��)E��͍��U��g������\^\�y�/u	�}������ܮ�C^w����t��g�Iʡ����W�CI�dZ��(5���cM�:��XCU��.�,��ج�YSW�W殌��\]�l�zs�c�s �%v�yȱ�yi���mj<��BZZ�V�	�Z����QK�4����q�Y��E�M^�X��tv'��=!!�K���C	o%Y��!���S[�����z�a��<������e�Q�;�ime,a�Z�j����AZ�h���(�xO\�'���^9���)�}�FJQbE�S�Y�o�X#ji�nl���o���n������󪫧v��<|��o8��:���DE�E�+:�~���t���y+s����k�^u�р�\��]��3g�n*}�z���ʭg�����۞�Z��z�F.CY���u�Ë�-��y˴��n�֏�����f���W�)&��!�$�DQ�d��c܂
�f4K�e����m"[�@D%���3L`�/Lq����ċwѦSU����Tc_}�(��m�X���6�h������
���9.���$�#���ˏǏ�Ms�P�zw}�M��������7��1� cȔG���_
�G�RYߍ��W�P���zU�:Um�櫝�����r���V�2��)+S��FE��}T��b�����G۱8jڬ�^�tc��a��H��m*�t�Y�iOLh��@wI$bh�p�9#�73�o��٬�w<N5d"c]tGF��i�����G�Q��Ί�蠒�k*�u̔O\��d��a��^�k׌��w��˅wôu��.,/�/�_���[k����g\x���ɯw�:+Q��;����k*w.Y�1ZX���c;$����;TJW���OB	L%=���|9�w�}�ֲ������:fM��q-�--��h�(�G"œ�<�Z�(_�+��4�aJѓ �B�z����O���lh�
P��=sw]�ۈM�ш���l3,��h[��R$��6�@ؘac��B�J��Ɗ�Mp����5`�Ru��9�@�TԘ�	�J����|�kB3�
���bڠ����F����-Lv�6��[��Y��lߩ뎚C���oΗz�����K�i���a�'��0�*��q���/��̮9�:�&��~LZwl��b��x��uM���\�zwe�[Q�[��=������/�W^�
|���L+��c���t���:�7k+�QYTtN��!���T#%�~i�$K�>�$��G%��e�ݚqk�8��xt�CJ�ݪ;��SH��ݿn?5&���C.�����g����^Bk{ȇͨ�VEV#a1f���T��F�q���jґt�����ru�{�g�y`y���e�}����h����5M[Zw{vV^T��5�=J�xW�:\h�l3
���_Y�]�t�ͅfX�i�x�I6��!���V�9��ݥ����[��h�%�����-�#�5��\�����v1�y�L��i�a�]�d�81.��	Cy����D^��i��b�d�KCI����]��Ba��`�.�xm�*������r��Na��rK���66457���,���1��KοfΜ���ȟ��h��e=߼�#7����P�}�G/�`��O���|�c�v|r�����m��O�n_=ؒSY��o���n{�cF۷V_�@������<����7+��{Ǩ��L�^2�ȋr��i�iR��%�6�R^2]��6Z	�.�rO�ʖU���^&�ԅ�G�(GB���K��D]Q��آY�-��آ�b��-j(�����
�b4Y�0g<{stȷ�w�o�'���3��/��|��|��|L|��s1���Vn��2�m4^WG]à��_jtD��#��SG������GMge���J�R������Ӭ+�R1�R[������4��7'��L�Qq��Vo���E+�������VN��6ֹ�s+�]ݵd�x���6���}�e�a_U��������5s�؛���;.3��u��zS]q������+��K}ld?�Ɂ�t��-�&�R�1�$�x�h�t�c�.J�T11S�q��˩'Ͽ�����o�ԏo��|��	,d�>�$�mf�CZ#a���&j�����Yi�H����抑0a��l�B��翑Ӧ&�˫�Ҁc5 ���*Jf0�|�.��f�0f�;�z��dt��G\#�5����2X�����U�+ɋ#K�E�k"&�n�L,���RR.t�|�%�/��D��PcIZ��BDL����nE����ۮ�}�&;m}}nfY��[�� �ݷ�5�722�����;>�%��aKV4�����g�ԓ�񌅼�y�ὣ��W�ԋ�~;An��	��v�,�  Wa;Q��6�'�6�4��zf�6	rn�*�L�s���Ý�:ݷ.a1�gf�M�y���b�F�L����)�'Â��1��k��@��kB�J2�"].�&�u:1e�����hy��B��9T����4�x\�>B��jnà*���&u<ȡuL��~�;(ج�Uߺf�8�]��ז_w�/.Z|�7�����n�,������sj�ۛ׌����uVM�;�h��G���_i*��
w3�橍�R#͍�j�K�(�"(V���5���N;��3�{�W�^0�Whĉz�2�l�1�
�tN�QMe�s}��k�b9��8��"R� ��8:k<�@�3�[�n�9�7�BxZ~85�95�D
�7���7����M���"��M�m�6��r�p�<d1�tF+&a"�LS+�ݖ�Vq����W��ʥFi��\:O2I���d��EbR��(3]�36EH�%#��!��ʦ?'�L �;:�^6x��A*H�x[g�Mgދ��np8K���֐zk��$[�(U��9�r��ܷ�n&�2��$�Kl�z1��\=��o�Z��6EsJH߅��]J:�2�aJ G�	�'����7�A(!Q����v���q�dɑ�S7�[��>�q�ނ����|���YV�	v���2�L]�%�-�Zӥ�v��I@	�RJ�Y�2�<ү�&C��F$EXIV(Q�n���Z`�ۊǂ���H$U!��FJ)�LF@΄Zf�=MY�)"zs�n4��z�:X����;f蜱��������ķBǜ�E)V�hR��`B�d<B2ZQʴ"5dH��`�}��˄V�jDMp�����J���}��4�9������Z�]/�<3z��9"Ko��~g��U�t�ԉ�E'�	k��ީ�
�8�;78w嫁�_lM&s^�E4��	Zܝ�_7��>`#|w3hM�>u�>��1F��@�%�`�z����k6g���JyiV����+�l��<��(�Pn=DM�����ǰ����@�m2[���Ự����a%�d� %.uvM_��׿s����s����Ʀ�}�������2ɵ�������pem�]taq88zǔ���:��<����]]ή�B��L��d!��]Iz��瑭�K�%�˽N�����e
6I*?� �5("Ȫ{|\d�v�P��Yp�N�J�r�Ά3vٷ���v���@�'Y�" � � ze�dZ$kY����q�|�`>�=c=�"t�Ie�6@���d��ѼG�%=.�l��Q�9�1���Q2�t���.��7�+{�>�g�g����n���Zv�+����KFS����u7_|�o�m37D����(LT��jQ�R��g�'�����{��V��ޔ�8e��e�o�ʟW<k�J����\��"����֜A�Ƽ���+7���Ͽ̱�L(����f���pa���B����!(l��̘nm��*
����Iz�,�`a�W����U�ѽ������{үd��j,�b�6W���6&������RM�p��1�"Sf�x(�MW]��l\�(HR��ɻ�\��]C�/���O���>���~}��A�g��gu�N���f�E�{�$���O����L7�{*�NSKu�e��}_�fisK~���������ކ�0���h��qk-��56dG��q������Ǻ�.��;=�]v/�,Q]O����wk�s��l���5�ھ�9ɹ?u־�zç�z�B�`�wF]�U���ou�'g���5CAwܓ��sn�6s6��L�����c���b�s`bf����7w�i�>�xp/��)I�B��.��l/�ͷ���o�hX����::jpcz꾧�!������9��fA^e�
�\��������I;��X�6�f�O/����h�u�5��k��<5���Ҿ�6R���u�&�`�&GS����RE�}�z�d��7} -��sOtr��_O�w�W`�6ɭօ�B�\k�У��n�ϳZU�$K�"��X-V������IDY�%�����l�D�+���f�&�=�{�E�s�~��#���d&`2��B�iڬ��P�j�H��&����,��;P��bIY��
�q�
��n�ؕ/	R�$Ht��< t�^����/��
�~=�G�{{��؞2t��:�/%}'��V�ևM+���������~�c�}�<5��< [����~_�����]¼�"*���=&]��Ƒ~����Z2!�������i��/x�c�G��Z������.��&�O�7�׶��+z,��-9��l�Y�\!@9��ՒefN��cil
C�pzE���9]ʖ,��kjji6l�ة �L�\Z~ 5��@��9#�'��C#.:pwiC��I<A��&��$Y�[�2����ؔ&*��;�h��{��9N'U�f2=L�'�fo�s�W��
�:����w���y��HM���磚��I���)؈�B���&c���m-���p�A�')���P�I�%�ݦP ����^`<��@���){�n�Cͺ7�3S���~h���~f��kjk��$�J��d� }ۊ����A�es,3s�x'�ט��2�V�=*l����`gSq���M�T�;&��y�}���ͽ׵���-�ڝ�jZ��\_(+.��<3�cm��nn��v7�!M�/ǿfE��E��`~C�z�߬�G�⎳s��)%�:��՟�2*Q����sR��E�- ��Koң�!)��TS�%鲀�p����į��e���u8��C��Åy�T�?�W��2:��|b<�9U�/\����q��F�����ښ�u�֥�hA�ׄ�����TRokr, �.Gw����M���}�=k��3Ko%s��ٙ�su�R���#�vK�K�=k�Վ~�&Ŗn��0�4䘰�h��d�;�-��	�� ���>�FR�0��]P���4̖��n���J�W���ƛ�,�A��*�+�f"�&�gu;GR1��.ۻ�k�9t\w��޼�G�m�csn��_u��rn��X��{ulUi��},�|�a�WNK�$~F����YRӔp�����n��
"њ�-h�����,�x��(�T
�|���-�>�dAQ��&�-�݋ү�� N�yZ�O�����;-PZH�z��(�p������7��H����p�4�V�h�H�=a74c�֔���U�F<)�����hU�H��EM�$�&4J��/b�G	�)���	����6ֈ	F�	l�^:@p9m��AV9(h�ֆ	FtgOWM�{����f��1�"̺h��k�⎎�n_��N���j������ލ�oKZ��,̙;�7_���y�7=��{���}O/l{�^bv8�F�����(%?�j[o�XP�~ovx%���/-x��m^���%F��d,!eS�v��K�q�L��r8ʦ��r�^8�L+���]Oۿ�LS ��HC���őYE�曂�b��i��6Ӟ��IVT�
�����c�W���ʢ�tD��9�p���H��I����`��`����	|�|���l�[��("��;ygҷ��T5K�7���X�mw��Β�c��xYw몯65�-�~ǚ廻���m��n��5�taI�7Ƿp���>}�K�-+�B^x������S'~�p�&%/J �B��F���os8�d�"E�H^�;[ l7<w�K��n��ʄjڤE3U�q$21�̈Lm���P_��Ɍ(VUfd�ȸ���FZ}�1�hssJ�U�g������풩$��@��	T�uȉ�߃�<9��}�F%�,IO7}��� }�M6�ѩ��!h��A�=�q`Kn^@&0�Ť�-.�^�^E�C��|9��>�n�K�3�3Q�"L�bE&l"0�	��O�|W��M�1����Iq�ˉkB(u�x� ��R2}��1�'('ݷ�#�v����^}B�PJ9�YK�����6�)|i�-mm�So�c�%5�����)ͽ7
��覅��+*� �">�&�m��On��/�s���)V�K���J+*���͡�8�+���h�z�j�,�*dR.%Kq@m�Y`���I&��d��<їIƨ��u�;a�)�}��"��0Y�D���xƵ6V�ճ��Z]#�N3����Z�t��lW�+j��z��s8����zt/ �zw�Uݥpv�v���=�� �-m�`��n#���� ��J��̇W�5�L.*�5�ՙ�3��t���C�"��E22a2a2a2a2aeG�2�O�{��.Q��i�Ӊeư>���)� �I���\)@��r ��L�3a�z�1�:K����P�T
�l�w�%��SŲٗL��W\;﫣���O4�4�siQ$������Y��_}ΕI뾷�K�7�$�E�?��cKՐ��./�Z��N��'�=����T��cos�S��j �M���d$K�V�ڑ#9Q�*Z���[�<2�H����fY�4�HH��e3��3��]�U��J��y�qWڐRj9���Z�&�D_�o�Ot����U�-_��F�4Q���[I;�k{6o@���o5[���m�Ř��$�ݰ-�5�*YɬS6���˓�v�_0�3���`��n��4SK���F�io�3���ں8�˞�v��`��v=2s���3��\���1�Ͽt��/�9vl����uTؽ課��m��A'�Ă%O��ҕ(+����%-.f�2�H��ę���=�h�4v�d$D#�a6%+�&g���4yO��,�RDA&�D�`�,R��"�*jz<\a�w�$�3M���F���Yen��-/�����4q�
Ν���c	�}LN�5Y�y� �{:��v��6��uY�92������
�!������*:�.j/��J�&DD�BD�X[����l��e-j?�ɋ^-#�g ��(�A��4�Ħ�Qd�c��d�c���������R�	V�'K'8DA�J�E6"�V��w�	 ]���;z[_�
2]�1Z��\,kE���t�,�mY:�4N<NU���Q�ʄ'�o̢��I��W���R��Lk0r��l��TڜSY(��eAD/�
���`��U��]Xb�����N����(X�G��n�5������ޭK����X2k"�5�|�-�j���ز@m��]�#����oy��F�裡���48���֧33�Z_���ҿ����9��X��;V�xOm'O�U�k\��w.��Բ�;��~`���n��}��~4�|w�����J[9���~��v��2��?B�?dI6:G�)}ڤW{v�`�~����n��Ϫ�볤?�0j)�5uL��N��R��S��X�Cl.F���`��L�&�@��5�-��
}:�} �d���Z'�3�^���+��D��1zA�]J�.bؘ� �4�Id����.�:��1KKC���8"��VQÆrL���|��Ҋְ�R<%Ph�혂/.�3�V��J�/��*�zUA`Q����o�����Ի����5�7X���`G�`��*�T���8YIN���GH�V.:�F!�Lo���2zA���&��:��}��d%}D�EvC�����n ��q^�L9e��&���F�i�{#{�R��Xpwk����ꃶѶ	�f/cq����p�jT������6�]'�|��=�e�ݶ����W�!�1�����c����_.[�5swVV�
�\���9��Dd4�-�v��o���WnZ�����ƋF��������E��ŷ��������2zHd��H�D�݁�X���_�����~j�'T�)4;���p%��/����E���}�%����/�����(	V���e��.��v�d������3}tg�ec�#Ɉ��6�UؐVa�%O�҈��ޭ�P���"}Mki���l@;���j�N�]����]��j�5��&��'~ltJ�������C�.��Lo듯.M��	�ψ�[�a{  c�1�j�.%ݞ�¤�Բ��e#���V��&�1{ג3�=���mfg��Y}�?�X��a|�*��^��c#9�=O\?���������B�؋c'�t�"y�i쁱��z�ѧy�W������Cr�?bɬx��|�q�=b��KX�+��J�4���*[c�е0#�Z�m|2�X�e���]�&U_n�v�-�3͆�_j�q��边)�ͬo���`���iLS@f�����ڒ�r�Y�w=��%��6��>���;BI{+�4kP{�<���l��{t��ŗ�.�R�c��<���#^��3O�$�ݶj�H�3��<i4	mY�-��,�
 -�Q I�u�#n�����*+�R�4��^������KI��mi˂�2�9� �q���nf��W�ǳ�~�<�]��l��<%��%JM�&Skl���z󖇗$����'.v�?�D,7��˽��i�i~����W{�����į���~��EI����/F���u��Ep�=�=����e#���Z=:�������k��(��`6�����TVj�Z�Y�ы�E_f��*����5�OԸ4?$����l�7Ⱦgzh��DV__�C��g��ߘ���7{�q���=3����������#�~�q��1��+�X�C�$iɛ�Tsь���Xx^_��=;^�Q߱�e}{.��Ժ����BmE��Tr�|.CC�,�9�Q��n��:��֎���ʵ���v��hu]��}�W���!�+YR�d�~�lmVU�4�b����`n/ y`uY#V�j�l�5�'���]�^�����3�v�.�A�S	+QT�R�6l�h���:G�gK"�	����[�צ}p��tA���M�������U5�MҌA��5b�xs����F7��������&46M~���_y�1�r�6��^8��;��x~�?λ�����ѓ+V��b!�w�n���s⫨���U��+@�,M��6��~��![���	�	����{��g�-tX3#{}%��Y����$2�b�c^X�
�z�#����+�K�;r��2�ˮ�?�
;�;lxM�������g�Ǚˬ�S�t�,4>���wFC|X{b����fe�+�X�(�zAp��aCVXd@gB[&�l��X�vʙ)����>?�R��w���sn��њ��cv�����f۽pqMC��ۅ_�~����x�Y�b�[
���@!�ٗ�~���n�IJ�fN�٭��v�	_��ؿ�2MEeA�#�d����9IE��I)"_�ȲjBy$����y'���;A]y�b6{L�.b�-�>(
b��2�"�H�C�M�$�W���D�Gt��#�Z#�>�}�@��ĩ�Մ�Fݦʯ�DdK'D��K�J�=��;N?��c1=f:d�g�f�­zB�7�V}w��HIH}�|S�;��\��B �亍<ɸ�F��ͬo�Oe�n2ZC�n꞉�k�Y�?$�Q�[�M*�vQ���6�m�����ͪ��5k�n5��j��Ӭ�[0��&��'V4ƣ'���f��u���z:~��t���ZdAs⬧[�o�Q�d}�`M��l��3��k%�J�R�X�[�4yY �Cz�s�[`#�*H��u�y�r�u�p��Kީ^f�a��:D�8EmTbLAEV�B�����%�
��v�;���-z�����Z�n�����Z���e7�|�-�C1�AIȑ���^��;ƞ?�Sb�*q�!���R�uq-�X`��D|�d������M�?� �J��;WiUV+��K� J�Z��BW\��zM[L���A�ل�n����M��(a7�ʡT�2]Ht ����B�.Q�d�&
D����>�?��kV�f�4��	��6���D��ޗtvj���/>�Q�}�}D�9�	l�����v���H-����6�G�)�~*N÷k�%�T��_�<<~�L��Y��T��
��=Umpw�{��-�F���M��
w�;��l���$x,@��+D$�&�>�G�er���vD��̧U��ġ����n�g	��3�e���.Mz��t��>���}�W�����cZ/��q��`I�%=>_�%%%��X2�;	��D���n)*)G
ϙ�dl�O��b׵uu�7���]���{~:�WP�uѝK�j+�����*k��޹hkaArmr�&Ƶ;4�U!�ڐaʵ������Y�����[���-��/��*�����&[ű8��Y�	��b����޻�EUu����33�07f��a�aa@DTDDDTDEDDDA@EDB�������)���^2"4E2R3R#5��%E3C�����Q�}��y��{�?=Ϻ��^{��>3#fg|���;��W�ǹ�X!�=�P4�������6M���Lh��WefgJ$��=C�-�j�I��}7��j�gM�y�3ܰ]�zkU4����E�-o��/n�bM�!��󢌼�x�[�}E�~x�O���w�|�c��F"C�(�7��l���+�|a���h(�ơ��￼�jB'L��?{nPpv����TST��6<��l��L��&�w0�0+e2�.z�̜���yy��YrUL-��1)A�M��HH��cҍB�����1�����ﷵ�:�+����[ٷ=��}�YK �(_�ʎ��
?U���݈� LG�*8��hK���L�C�����������Sp�2a�GW��~&�5u��w���J�`�D���Z�>�a��7Q~~��8�)�?p�"�1ŀ� 5�ص��������^D�����$�fs m�
5� sW;`������C�{AG�z���RBƽ�GLH�h��-�'�<d�}4/#$7ק[�.��P������n��
ԡ$N�`���n���H�&ڀ��ۮ��������=�{�- �Z���ɽs!4yu�fo@j�FM�@�F�\�x��c�eB{��ݧcV����򎽽�ۧ>l��/%'��՜>�~�Z��̦�i�G�K7��ܜ镆�Z[���������U�t���t����2'���W�o1�1�^�J�t�R&Qw�8Խkg��˫��V��s�]��A�v��g4��p-��W�q�������3�x(E��W�]�������^ć�Z�ы��5�,�k����j4UK'3̏���k��mlmE�!����<U���{��]���M�M�i��^�#��=���U�jE�r��%�KjOM''�H�S��_K�&�T7���X�~����u���|����!}�x^</�ϋ����y�x^</�ϋ����y�x^<����������y�x^</���Ϟ;/�ϋ����҃�����Q�H�*�	67����Q�� �7?<����'��|��tE&໢p�#	���|8��6��� ��� 8�B�{���x�#	�!xt��	�B ����#��0�&aw��p��5�Û] G4���E<��G̏$��� �~4�	'<)Q/h�'���'����2�Q8Ժ�!R���a�ݛKG4?��wo~���㒃��m�W^i�����EC/�� Jr��# ��a��a��a���$e8INRb �p"��0�G@�H4��H�x�� �j�xts=�D�������>J�E	d�Iz"�y0n3��I$m&��I�9%�ځ�B�x�C����������oCҽ	oK�`�ہ=�@,O!���4�Џ8�Af���ye�H���Lx�E��m�m�̍�퐎�s�=�`zr�X�a�	/���=��*,�%�w�Bx�C9���^iQޑ̗�U�N��i�;���6],ʸZ�&R�:��@�.��Ә����E_"�tQ�\��4����d�����R�J��Pȿ��@�@�P*��ʔ0;�}̗ �3�v���?2#?�4M�r��t�t�k@�Hk�'C�dಐ���3��@�D4	�)hЙ�S����EC!�4)Ο�B�i�R,� s��d2���L�&�� �A�9=ZGnf@�Rw�V�4<�l(k�~�p��� �&A*Ν���:�XH�Lf����mP�)��S��.�ϑmg7S�e�N �m��,�68eY�4�v.�#���@��dR/�h���FJ��Z�]�l�F�R�@ҧ���ciYöy�|l'���t�B,� �P�,�ɘ���񘧐٥���4��3���H��d]&���<�f�q�@ɉ�N&�;��iz�\�Cx��+e�3��/.�KJO"9٨'�gy|�u�}��?���D2slOs�9��d~�D����q��M�o �C֙]��V[k)�Ӧa�H&��&+��es6�M�#���MV��;�k%���I��d�x��$�J!�hY5k{��j�֛�TJz���%�&r*ԙ �7g��C��z��c=��dmg=M ��Y:���t2��dG���i��:������g�Ύ�?խ���-Ml���d�&���g͠��������Lع��Z�u��s���_*d/��ܙ����ΪXo4���X~�K�wģmY͖vp�L��o�l��V����2��r����N���Wb9M�yd��j�t{��&��L�T����ֻ���o��H���B�iY�dH�Z�H<��˵9��{w�vp�ǘު����;��_�G�UQ-m\Z-:�صj��4�3�8�f�c[,��q�e�����ޜ]w�Ҹ�X�ŭ�7�w[��$b���n�g־������OMl��j��d�vְ�k���h�R2�;��d��r{v�>��+��"7�٬�x���������X�N:J%�&���yz��2��%�-�l/�m��Zto]k�����nW�3';���Բ���J"�dk��fa!��+4Zk���S�XҸ�5�u--�	���܊O';%�u-{��-��Z����,-#N{�n��,�����cKT�'�,N3i#H%�٦�(1�"����Of#@*�AK����7O�V������-�MG�ZcƳ�J�ZӉ�`�+�����o�sV5�U�Q.�&s;����?��X���CQH� zƐ���f o9q �Cj8�t�#���d�F��	�F�xǶ8����E ��4�GC[�nO���� %cH�C 5
h���RF������EC-�F3����Hc!��:���Hzl��b��H.�/�=���Ǐ�� |t�8#���%:�-�6������SG�F����9���&s��|v.��p�>�\�rX?q\^#<>�6�mV}�"�h����0�>� ��v$y�Nf:�h�?�3<�("�͊]�~d6X�X��Ъ��ٱ�X��^w�H~[)v~}9܏hn(����G�X�V8כ[�2�^GK�OJ�%3�j!�z�ѷX'��P����ᵵK�U�f������V�i�`��%:������Zf�g�{�d'Z�K�=MZ��6i��̐w3<=Ϗ7�7��p(����Y�5�*��3��оP>��-�m�C�_s*@��G!�3d!�!>b�o)I�ȯY\�U��]��.�v^#�!�l���� �U�����v~g	Ck�Ȝ,vP<��;M�JG����-Rt��:L���AN#�5?f7��xʤ`��'v����1��RD��hb��*s����)�Vt�!�U.��6c�2�Cfq�h)>�k&3�'P�#G�)�X�UG%O�49kb�,?�Y�m61i�S�e����:�"T8�<!g��i鹆~�r���$�N�nfW��(4m�����u��<5�0�__�^-�4�0w���-��_�A�y�����Df!ηW0}����h��J��~��'���G�7��3ܿk`�����v��=�ϯ�ٝ�����3s�4se�T0�GL%E�.�(
m�Z&J�v��N�i����?�w݈��}R������W�C��X2=f��9��KVz�fޝ%]�uYpƸ͚�c�τ��1s���?)�_�w�¬wl����]���klӦ�,�qs_���O?��rq���!�-o����	�$�o.��[�{hrE��|�hv-�����K��k��}���G��W&D]�c������G��'��6���Rڰa|���y�&?x����K>��n��E�'������4�~�����=������'Hz!��Z�Zq�q�4���4�7��J]$<O9}�z�����n{�^��|��7�[�	���4fU��=�љ��l�пf���s١n���X\��7�<�<�t@i���&��f�������3�e�|&L��=e2N��Ι�:cB�t��eīH�������/��?D�E��#[d3�0��`֬Y�� -�oZ�5+�x;�	rM2�V���Vy�H��c�	�#���fqr�%i��w�X�ׇNg�W�����~#�Tp�U�d�)c�O%����TN�*Y�؉����B��G�4|'>1���7�2����6�ڟ��-|����}�p n�*��B��+l�k]M{.�1/��:�6��������0c��o��j:��_���a���_�</�|9�V�x���Ƌ=�||����><��kY�?S{�*:�|���O���}���N���kgHڟon����Y�	{���x����vt^�L^�q��w�W��%�?��Y��\ ����j�Ū]�(o��_����Ԛ=x�y�_�i�`7��e~j�a��Y�*�c�?%g�����o�'�ufm�9��2>.�yN�?z����C6o���ql�ߘS���ვ���}pt�"ߞ]}���~<�#��Ӽ��J�H�o_���_<�{���Y��M��UG�5O�����T8.��(�v>(;vZ����ۙ����=�љ��1}�j��o~Q����[�-�~��b.��Ĺw~�����������뎔�_~�`�u�t>�W��߾�������)G_���{Q6<���&2��n�F���]Ss=����J��K7_]�>Xwd�����˻�t��Teڀv�q䵬Nc��	�ʿ�E����o��˺��ݴ�([�u�2��h]ʂ�����<�*�D��>;�Xe���<�E������lh�:,�/��E���W��Ͽ� s@J���.=R��w��5пK*D��d�n�ڹ�Ȭ�k��'���w7~:uˑ���gz�i�Ӊs;+��;�.��]�A�&[���f8�X�����A���.r�"<pE5�h3���LM!����QU�j܇n>��[��|�����wkD������_n|o̊qA���K�V�o������v��w�G������٭�-х�?ڤ��b����\�v|�CѺO�Gdߞ.�}���c�ۦ��߼�Qw5�eQ�O�(f����J�۳�wX�X�N�%5.>�.�R��!�*����k!�!��r_ԴS���k��ÿ��7�GF񖍅S�=��^�����c)��?��X�j��Y?��Zs����ߏۗ]�x�k��jhz���C�+�z+�R~t`�;��4��|��셵�x����_�Z7�T8��G_�G{�b�5�ɚw�t�4n��}������6������v~1���2���zs�_�~���hL�fj������򃊗�+�ۘT> �۝��j?�?|CR7u�6~X��-�s����_O|#�����k��6����[;����g��k�̚}��M���]�+�;�S_<(:��^~5t����O�1����Px{b��}�ux�wRm}@�;.��f�ܩ>�e=�^�睟��l �a��0Y5)��~��	vq�B���޽�J9��F?'��]�]���vf����o�L��Lwr��	ɹi��3r'M˙�;;wsws�������������Ռ���#�?��u�3w^�)r���)>N��]���{�݇}|�gM�Iz�����8�lp�������Ö�X�h�8���xy_�"�ު�����jz��{uލ/�R�r���tq������M���,����͙�N���\Ĉ����<#|:n_8td��*��WƲe�7�6��x^���7�V�{tBq���Sc��_�.��бS���WO
����(�
�-�5rvU�2��u$3G���{��]b�}����oֱ�z����d�S���?V�6��?Te�o���@#����of�X��g�.��v��x`�2�)����W��y�2������C�:���A��uI8b���Oؘ�_7�ٜ�U��n�8jz|���'�<�
��J���]��_?�f�@�ؕ��k"��p����<������aеl��C�Lx�Ͽ��x�O��B���}i�T�b���/�]�sJ�a�Ԕ�Q��h�b�{?�^��'�%�K.���_̾�fm}/����o�5oE^�;���ۖ_�孌�^/�'�}���/�1����Wg��#���rv�&���S�9+���X3��W�%7S��V�i�s�F���1�A3�zwα���ݻ�u��B�0y���տE���W�:'}��o��؇�|jD��m�/f�%���B���Y���������˟�/<6<����E��{D�z8�˭���Nw6�� ��M���~�k�]��������kֿ�镍[r��G����c�}p̒�"�)+w�.2�f]Xs�������a�$m�Z�[m�_;��EC�1�S���<�"M�n���|�������o~�\���n_�.8�1v�Όދ��Lޓ�^��˭�ʧ=Y쟹����%�ߤ�{��y*ݻ�'��.��v�Ӳ#�̎���3l{Q٦��v��ОY��b����mV�%�,����[�o��ߔ�x�*m�"�Wj&�\Ϻ����~��%_�I<=�y��Ǿk���TM�F��s�M�����
$�N�P�X_��W\����n�N�ʆl��A��7w���@"�����~c)���4�4��s��>Α�|>>���@6$����x�ua�^S~M��\���x��H�s�)����U�'(�����;�H<'��yE�M������II'.��K�}�3uޑg�ɏţ����M�y�?�C���6�a���l��jfƶI��N��3q��!��bP����n�7�N�v9��+�m�?$��4��/����Y��z���J���8�y9�=?�t�֭~�v��]//t>�s����.��[�;��^]vt��곐&�����;w}�<hމ��Dǽ�֭áY����X#���}�ц
f�[��[�咢7*��v���{��gP�U=~7w��:�?J�Ov͸�9��q��;�=�68$���Q}L��������~%{�txĬݏХ��t���8���|j��_z����>�RS>��Ճ�r�.��b��e�{_ݩҍ�鵷�4�m��1�>i��,�����_�Uwk�/;}�����+�/N�=n��G�I�r���﷦�|�����C^z=|Q�]�W�6���]�G֣نxo���+JB�v]p��P}~mtCqYeDi��
����[;}F�k�ϼ�8�VP�<�^�F�~������SA��Ɠӥ'���J~���~����� s��ԡ�CJ/�o��}�6k�d���8�,�\�y�9�"̅�ka�o��5�_�o��_i�_d��N��|����}Z��)U��f�N�0f6yjrΜ	��}&�N5��6@��������[�q�36�3�9 M�>-Nk��������{7��;G�s�t�D�j�b�K��V�ʉ9�e���x�<:����ך���!<���}p�O�4v۴rlڂe��1l�i��'��u���ތ�-{2�J��O���{;o:��ˬ��M�&���<���W6/�}��t�W�b�?�Vߚ�x�ϊR�>^S�Np��������k޾��|c��}��du�q퓎�j�/��=ϕ��Hz�߳]T�z�_s��W]��Y�g`�aa��w\�u�'������_�}ugC�G�{&��5zѤ�i~�{(�/�Lyy��QI�?�{ȃKo�����J�g^�J���ؘ���\&�\x���G�T�K:^�v����c'��2�f�!�Y��;g�*�''z��ag��}��x�>��[������Өn}ľ��Wn�){/ߵu�j��M}���w;|bÆuyy�Ǒ+\��5�=���G_N�l��˿͘������9���u��'͸����7�Ͽ9��'��[���.̘:��߿=���Q�����������זc�\_�z�Kqё��}�z�a~�'s��7uj�71��a�������4E����\�~���H��j�|8#�c�D���(�${?��2����V����\�;�D��~��{o����K`N��"�3ǖz�{>�+�O}!r�G��;;vN���9�ٓ��b3��B򶹸�6�|��˓�����y��3GP��Cvռ�o�q'}����u%���t�d�����,�֯�o�>�]Z����x����Ԙ�OPL^����s\�vq�����_ސ�{��?�/N����w�:ua���Q��K�.j*�S��0���c��|>�>�����g<�5����x�l��z��K�sW�O�(LE!��{>���p�B����M^r߮�'֞t�?5�4�{q�ʯg~����~�X��m�_�"*|�$��,7�i�~�"r2�t}�	�S�	�
hGHr ����"���,lr�Yci��mR�yk�OJ^������߭��S�ւ�O�_�_Q��P���q�{�[]�����~'a���ov�T]���3�Z�ߐ��p��������
iީ��3#�Q椲E�+�?�n�A]�!Y������:έ-�S���`M�\��=�Wl��q���طf��u�ggbU�_IJ�zv�.8�vŜ>s�U?��0B5����N,����v�m�M���st�+GU���'fi�)�7�?�q���AO�Z��w4�WF��wm�v����A�_��8y��e��ƊA�%ݝ���=J���WTwF�}��'7e�x�t���+���~R���=��|�聈�щ����K��~�����j���k��^�:�.���g�2"D1bF�Ɓq ^�ȁW0N�k-��L����G1y��̼�\f�2�"��g��4���(^W^W��x�O���K~"o*�Y�����<ޛ�/���y%<3o5o�y�����!�[xG�?�;
�1�E�/� �w�;���7�`��?�Ŀ�(�U������7~���ȇ������lV�\C��u����i�C�]?�H������v����s�+�����/����]3��Hh�h���x;��r�x�p�������>A���a6�/	_����/n��m�m��]�	�eB�������a}��� �~�=��>�>���Y�O����_�_�b�� }��������=�K��_*JF�(E��Q��}�׊�!ZT*� �Q5�%�(q�xbĉ�DD�ǊwA�n��W���_\���g��I���$zDI\%=#�)�hI�$�ޒPH�+	��$�����GH�+�|�$�)�L�J��%ɂ�I� Vr���"J���{�HO8G�C��8�8�w|�C
��3h��� ����`ģ��!�Ųv�� <�&�� ��%��m>�)C<��6;��m��6������w6' ��9�gl� ��`������˴�ds���"8�iYӣ�o�?.��'�'�z��x�K에u����RO�kD�*EW�� ���հF<2K!��O!~rNr
2L����fOJK�A3�s����IɓQ�!^D��5ڀFD�P�Șp����L�1���!<��62���r�x�"9��R]c��q([%
كL�b��"!�"��qb���'Aj����c%x+�U�%���PB�5{@p���#����:e����c�"��W	�'���F�iѫ?�P7��� ��D�����zi���\�`�҃�A۠a䄴���R]��憌��P�:"O�	y���uA>ȗ�A6 v0V{X?1�ճ�(l!�7�%��J��螦r���([JCyRQT"�Iͥ�Pk��T%u�:G�S������t0��D:��K/����m�*?��O� A�`��C;�����.�.�.�.�n�]��9�P�z	ㅓ�[����1������(Q�h��D�UT!:":+�)z,��b/qO� q�8C�'^,.oW���ϊo�K����� Ix�<�bI�d��Br��M�c�P��zI{JI��<�bi�t��BzDzVzS�X&�ie^���A�Y�,O�XV"�*����Ev��X��ZHj%�"2+��5%��ћ��ʹ��ѱ�B�|�D��'��P2j�30���T�^W�^N��g/k/�崗_^��yQ��P�xJ�!;���6�}��dǷ������G��u�����օ���#�i�X��#,�DҾ�O�u���P�>�`K����L�V�t���րA(š$�Ve��hZ���b�mF;�^�F�Q:����\m/��p4������]����V��r4��X�G�Q.}�ާ�>�f�)����r�{���3n���s�K˵d�F4Š�]���
�b���h+څ*P:�N���2����M	)9�����O��¨A7�rn�E,�<��7YZ�i����_s���YZ����s�[�}���Gp��ؗ,=�i� ���\������q��wȟ��YZ�ͣzK��rt9K�8Z�ү9?�uG���^{��-"��X��3��-ō�{�����9�;!�h,G7r���'9�:����xz?��q4���H{�7A,
@�(N(�(�"�Oq�:ŭ��8Z��:�\7����V�t(G�U9#{֞=��e,=˭��ͤt/4-@KPZ�6��h�D��:�Ρ��5�F�G�(%��L�7@S��b!��B\˅ȶ b[D����@���w
��U�s�x��L� ���>���D���4~�*K����_�V�"�b��Xz�[�+4Go��j-K�q�];���X���~��׍�,��k����܎�m1K�9�����g�����ͭ�mnw�}w7���Y�;g����{�Xz�_�GO������Cn�p�y�Q�/����ǜ-<>�ҿ�r�K9K{���'�Y�ĵ�t���E��(�?Eq�th�}K����[��d%g[Ʌ�"7�_�^Ե/oS�>�V��Τl�9���v	�� �hZ��^pz��������VA	���g�3J��r��Z�q��l?����<�5�QkQ�8���kX����1�����Z���hG�H|8�j�͝�K_��
��q�K��gדj9���fqt�s�s�ӣ�GYۣd��Oƭ����,��39����6p� G�s���ZR�j]�8:��]���k8Z��sm|Vi���>��h�3K�s����<�-,�#+��!��ɛ�˪���vP{���^�EYɻ������as{�mX{ٸ���nk%״�;X��8�^��~?v��^�
��K���jl/{WX����Rj%o���Z�eV�^+��J�������Vr��|�J>f%�Z�uV�9+���|�J�i%ߵ�Zɍ�e�J�Y�B+Yf%��d��l��=�do+��J��{Z��Vr��j%�Y��Vr��i%�����h+y��g%'Z�)��KME�����=<"o�m��v;�]H�uK�[n��.R���@�䝶���.��������6���:�7����m7�7yC&q��P?IgI4����'oVG�w�	�m��}���0D3JF�FŨ�qb����1:d��3��+����Lre�0OлL3ӌ�x[x[�
�1�yTL��D��o��)�Q�����`��n7��~�}��}��hj�}�HL},�#�E;�7��H����*�Zr�^)9&9C��~#��?r0;�w�7��wh2B� p�5 }���-�{�X � �L ^ f�@�`�0�H�h�X��� ��F&��� �  ,X�A1�r�@�- ;  �+�Btz��i�� p��
:?hDHB�uH$@� Z ��7�?@ �"��p�W�p_�dP;��x$f�W���
$q��H�����Q��Mi��ZQ��Ft\tJtVtQt]T/�'z$j�JT/扅b��P�ub��S�#����P���#�Qb@���xq��Ð
�28Ȇ����q!�J�h�X%:+N� .��7C;ۡ\6���9�J�\	��x�a7U�� �Bz-�׉.������~�8an1�2@��y�s�f����߀�a8��m#��cϓ�� Z�xQ��\��2��P^ ��$"���:����.J�X�hD��}�q>��#��'��,�|����$��9�/���ۢ?� �"8��x�λe��%��dt�r�uq��e�l�{ܷ$�!/�c��I��s%��hI�$��!�� /I�dJr��t�l�2�F2O\(Y �,���B)@h�M��N������m���2I���d�S�-�oY_�A�)��� >����J���do���Ж5}�<�N�t�C,��j�\:�j���i���в�-��U�~��%8�I=�[�1E8 ��g�� ��UI��ٲ�D � ~�Yq䟖��<(#����V[�(����]���}�y���I�- )-Va ���ʆbh�;\���|k~(���R[(o۶���E��b/�]<+��^[�p��]���������2�o؃�Z����|^��>g�OR�Ck�u�l���V�,6Bzy�O���ľ����I<��V_&9-�#նش�ߪ��lYb�xI=@�I��[�?ޟ � �Q2O�~��{\:��)kٲ|�%1��Z��-q�*����	� ����e�n��a�z-{Br��<���d�ă���=��dO<�F���,M��b��[� &�׉o��NȂ�v`_��.�Z�"�gmL�lt3���mI�@/!����6_��ئ�r��t	�uV���IZ|�t��Zq!�J��Fؤt+���/��"W�\r����S�gK�KOA�����$��������ҋ���0��xX�'�к.-�1�zܺH�{
tJ�+}e�pf���g�爽p1�j���:Gp�U�$9!�{��� 9{��zeB��$���	�$��s�KI40�����IZ|��S惡e��
n��Y �s�9��ږ�o;�zJ2�b!q�,�,J,Ā���]���}d���$��/ˀ1b _%�u�ͅr0>��zZ�$8w�sn���;����d�"%�(^&�^<`}�7�M�kp����@R�<�7R��FN�ؖo��tJ���N�3���7�t�g���P�"�����y􄷐�����<�K�eP��=���.~k�"�0⻐vR�d~�e�c~�<���[�܋�U�{�\�p\RA������"�����MA̳)<���[ �Pf?3�.�9�A�kÖٌ1��	���&2�#dJ�B=i�/��<j��������N>o��s�$��S)I-�ƨr���|� Ŗ���AZ��rY5��!<j
�<��y:�F�������H�����x��$�{� �l�m`n�1�\��jq��ȷ �1z�ˣ{�W7�����dT�����U����2��$���2Ix��b�r�����z����J�'��#H� _l��m1������r��7q�<�;��HIoNo�o ��n���c�1�22[�̚&<�5�jM�dل7�H�!�_��r�7��t'���.ǽ�$�#^e�@�7������I0���1�#[���3�B.�R����A�5x������r2�rVKxe��{�X�-�u?�OF���V�K��¯!s�%�ѓ`[��5��%'��`Ob��1ia+�/�6X���%�������b�fѡ7���d�kƹ�p.�/��xb9�dEM"��d���obi�6x�ד��$XIFU@�b-y6��X�~F댭�P�Q	X�?����G޼%�7o�ț����[2~3(܆����Q�@� `��e�7 n4 <�_� � �  =�	����� 0  �� �=��� �@.�Wf�- ; � T ���@�� 8p�*��z�!@#���H � Zl;�p_��Nn�3ޭ@1����	��_���
���|Ą?cLϨC�j+C-�V���.R_&���6=	{ zRs�v+�������x� ��������ݚ/�-^&~W\$�Ι'ŧ�?������g�)\y��Ӎ	d1��;�]�w�����O���������WZ[[)^%>�#�V%��Q�rq���?�� �����}Z $��G�[��M��}dG���@�W� �w��E*�p-�f��|_���g� b`��M [d2�f��P P����`3�v�] � ��{2`!xO�'s �'��ޓi��1������ʃU�������L��3 xPxPxP^@$�����݆x�A�n���� ������[ ���G�m!�Hm���x;����#��<=7vk�h�G����Yu0n�]Q(�F��������b��k��U�è�EW�m0U9��<� *���b�D*�ʦ
�"p���z���nbx�����(@[�ݠo3�~�y�*�q��O�gq>pG�Z�6�=@����+!����.���iz��!u�B�VR��K�;L/��b��|�_\6���K�+ 6⑖��:�D�� ���U�5�q<*(���A���t
���0>9��(L�*ZG�Ӟ�� mI�i[z+�D4��j�Ki!p���GM]�nҶ�C�/��IgS��L��:N�����\��.���ET%U)�t�3!���J���:��~(�A�%����N�6y��_��Wy)�� Xf� pM3h}o�[�S�\���BR���M:�;�Z6E�����7� �����x�U�5�����	p]�8�u�bD�o��~o�����T��]<f�B�{�pO��ۅ�q\�f�k��gǧ����lF�|�b�j-�'�_4���/q�$ˁ��ΌT�oA�������D4-D�Hf 3����2�
�d��î���߀8VϿſͿ�c��b����G���l������ ��ǉG��ţ!�})> >1� 1J�%$��ۼ%>_�Y�/�*	�t�Iz@�;�m�C��H�8�x��	c�:$Ạ����1�'���J�i<�� ���O�pr��i9 �z�i�b��$���������`	�r�U k6r���|D����8p
�,�E�� � � �,;A@�@���0x�  ��� 뼈���ј���H��xu	��������i�聟8�)�$:�Υ� �,�����U�6B4(��}�2^2BF�bt���d|� �'�D0QL�$���=L���d�2L!���pfj!,c�9*�����H�c��{������o�=��9o]��pd`Oj�?���Cj<��B`�s��=�II���B��P�����lp_����O�Ԁi�q-�{3I��	�������u�;$��\O�Ax<��;ƶdv�$��z�~/cڒ���.�
���l�!�f/�
Ilp�s$|��`l	x.���|�'��&�+D��1�A�����ْ���0ZGjْ�*���@�?��2L�O$��C�J�R�H����TXMߧ�NĿ�o@�C��'�ǈ��?I�$&�����K�E�'	�t�~�0
j(���eY5��(�(p>FpcC�(�(�(pZF�������-�%��(�읃f�yh�b��5h��w�=���F�Z�~�y�=���+΢Ym|Rb�B��6�.M��6�mr��M}~�`6e5�}�q#Y�fI�$������`���J�I4Y�$�P���G#1x�!�n�7�<��6;���VG~y�F~yk��lԗ����U� �Q�	k��~	J$�j'�U�	�b2��p4N%)h>
@���ݽ�F�NףQ���h4�OJ@��ǁ@��"��^B��z4=D������T��Q��kh7�&�ݧ#��/z,=5�3�<��_�);��C)1x剔��̡y]x>�3� ��r8	���@'p��_�� @Н�*�)HuD	&RقY�A��]j�`�`'���C[Oj���mꄭ��/u�6�6���v���m����wl��F��Ŵ�v�m�a[i���YN˄;�ׄ{��ӯۿj_H�)�����R�v�ZtXt��O�>!�A�}FtZt�>+�*�
Q!!�9D��6-�۴n�r�I��&� E+�*D�L���д�$Mϖ!`�"@)̈VrL ��·A@�UZ4@�3��Z@�SyH���	n�tv, �y��ʳc�l��p�W��_1���  ,&�h�?H��u�l�,�2�_1k8�@�Vl�����V.�+�Z�A�!���˃�!�p� �0y�<Q�"�$ς�\Hϓ��ʗȗ�WA�Z�F�Vy�|��R^%k��姠�Y(�-��S�ס�z��A���O�7)x���Y
���B�P�)�
O��<E �=�P��(E�"^��HUd(�3s�BHOR,U)J��͊�]�r�~y���Q�*���7 �6Ii���J�(EJ�R�إ�+MJ/�fe�2X�_��T�)�����xe�2S�T��(Q�V�S.P.V.S�����e�� �G�<�1֛��֘��|��*֤��_!S�U>T$��FE�#�1�s)��G����	Ƽ�`GoG� �E`o�ᎃ s�Sj��J�����)���p�cI�mm���y��!w���厫�:nt��X�ױұʱ���)ǳ��˕��x�����96�x*�J�R�t�y*��Sy^���eTX*UO�C	Ap�*F�J��8��$U�*U���l�����ᙪ��:U���Y�*R��JU�U�U�T���~��j̺BuDUթ�)�U�U7����Fa���ԩ��Z �U��r��F�W�T����ڬTƪ��u�<H��Vp�\��N� kt�Q=r��Q�c�Tg�s�	�ZE�<N���-W�⽣���T�@��5�^����/�RD����u�5��oQ��<Iߢ�|�a�����R�����>�W�s���Ҥ>�>/�R_U�C����r�]�CGHoT�4��V��w�ڬ��h���x�)�C;�-��L�XcP�h<,xo�yE��_+ߨ	>J�	~��Z�0M�:V��I�L�dir5y���S`�DK��XK�%��ׄ+�4��D�*(S�YK4 ��lļf��1�eث����ż��q�U��c��~��~<�-��S��0�����U�#x/h�k�1���e�#M��Iqĉ�Q:	�;ɜTN:'�������)@q۩�S��$E�S��
�(E�S����}�S�%��k�ꘫ49e`F<���|�S����բy�S��N��4�M�Ns11@;-�J�B�<�T���ԩȩĩT���i��X��K�T��2:���+�J��ds��Մ?�T�ka/�T�T�tN��tY-��o�^�n��]�Ԡ(��aǋN��J-�>
l��^� [��V�X+R��v�\Q����ނ=��|�V�}�ք����X�|��X���U~V�9�����`����a�H��s�c�x��1����s��L׀���ʃ`�E�a�i�8��h�\����lE�vD�&�V�#�v�q�ńh����bE�v��kk7 ��_�e`_c~����p�	1+N{@{�=f9�	+��qT��Ղ�h�jo�5ڻ؆����Ҵ���F�)E�3�`�ζ-���c�)���n�+j�b���j�^�~霵�2g�f��z�c{�
�%�|!�iM�g������9�h�C,���9�A��p�v�sNT
�S?	�J͝�p�t��,�1�9�9_���]���;K��p�1����6q���8�9�Ԟp^"�r^�Jm~-���*����]�\�y�,�\)oRmw�r��\�OZ���ǡM898�r>�LP�v�h�/ʛ�i��P�8�v�s��=e&��l3Ώ,��6[���	v�z����:�B�T��)ೊN�O:��^ç��t������(�x����ض�Ŷ�k�����'
]�%�Z�.JmRf�b����;�i��t��$]�*N5�Ϋ�ro]�n�"vS�n.��]�. N>��Bȭ��H��� ]����P�R�f�v�.m4�p��x�]�r�~]���R}j�8��j�n�=���6�n�nC_Gtp��/�=�s �k�^� (傜�Jt�.������E�bR�\��B�]��l���V�v	v	SO�D*R]��H���ĺ$���x�t�LEO�S�P�M��l�x�y.�).��|X����j���9��B;�.k\6�lq��ǥB�kX��9_���:�Q��à�$�c.'��K]Nkǻ�w��r���C�F=���K�J�Vo�{���� }�>\?H?L�Oԧ�'���I �%�����xBq���.�&�\pz��'.}��H���������Y�����U�ѯ����B��;7�D���b|�V#�T�ߨ�
1q�c�e�0�$�.u�~��R_���ןҟ�_�_�������9�����\y�By���9x/��"΍Ս-�pU���U�vbq5��Z��'����� '7k�x�i8��)E�PQ�
���ǚY�5�4��qL�U;^wU��F8��8[�B�����(x���<���+w�&���f�3���"^�뚭��:S��u��Ĺҵ v�����9E�k�"�y��RE�k�k	X{*�����R���h���E!��LE��.�kĸ�����|���Z�u�s�U�r��z���k��crݥ�;�A���e�Y�6�����K1�띊�ޏ�SO����ٙ�@E�!�5B�j3D�,3D㓭S�!֐�ۥU���LC�a�a�RdX�L�b��+M�e�b�����U���Pa8`8l8�6�p�0�P�N;� >�<�U�����>���Fî��>V���Sk�l�n�\7����<ܼ���q�eoFnAn!nᠥ�p�m8�\�6ȠQk���-i��|#��0v�2�-�-��n)n�ܲ�n�J�[��V�|E�����m���a�b�����\o�-w[�����ݶ�������U*bܪ�j`���ڵv���E��n�n��ȭ��3
�2�ʨ3���Fc���1�a�2����I�Tc�1�8S�1�5U3�Ku�"c��>!��1��E��NI��N:�v�.c�v����G���:�9�e��mc��;r�������]�w7a=�{a����݃�ø�-{�e�wU�J�����o��=�=�=�}�{�{�{��l�y���/s/v_��}��w�S��W�p?�~����iܯҌ�u?��u��z���p~p��G�~���a�H�o�Y4��B��[��܋M4>���go�x�L��td��}dR�}�I���p�q�i�*�lkغL�&��ɟ}#���@��᳖)�b
��y����M�L�Lq�DS�i�����&�����L��<v-L���B���j�����Vi+LkMM[�Le�7L{M��*S��[�h3�2�6a�rD5��"�I-�[ȷc���{�X�r��(D5/'�Yl�����Dz~�;��ώ�"x9Iѷ��%�_D�$�<(C��Q����(��%/��ǘ~ץg��ҳ�w4i*��R��wz�`.����Ϳ�$)�p�t&I��)�2����_ �")��@���}�UU��>�9��s�4�4"""ш#ሄ#�ӄ�H��&$$$BB����������#$M��#"���D#�8����}�s��O �����^{�}�^{����w�>� �)��S��2�8H)�)_��-*���8N1c��8�݈�f�g�g"�n®�<��i|������3�]������q��̹�	鍚+�eJ��x%�Lǚ�q7ʳAy.r�N��S���U6k�*G�d�Z��0���n��R 凜I�)@J6㘝�w)�3��ٺ��L_� �v�c�c�2��tk��q]�7���a6R� s������HcG���{��U�_���c["���[A1�!F��L�z1?�ģ�e��s�#�Y�O��S����7A��Єҏˏ���)�q��$o"�!
��56��&�lG�{�b��l�M�lu�q�(�ʻW٪[��	��|��G�@�����-�, �ΌI���~�G0���咶�]q�0�ك��|�����s#ǩ- r��;�_g-����u[��jg�nk[`-&�,d۰&�F��Ne�0 u��5�|-Ti�k&���{�_A��l[�{�[�=-b��9ƽ���ׄ]�MMC���[A-��CkhNu'��9����U��t�A�?�$��y��V��kx���[������9�u#�owW-\mw^&���p1��P���?s���s;���%R?0q�tG]lC}C��L��|��2ZV9s��橧������{��{8n�Gz�Z��ބ�����=M�li�SQ�T���tV�1���������1�����U�	��n�s������2h&_�w�a�P�2�6��{�R�9�,�����<��6�Z1ے���z`��l��h���C�S�<J��r]X����
�I9�e��ڮ�q��w1�t
�e�S5��l�lu��v�~f�;�`������v��\��>ƚVQ��-��ߠ��m��)���@3�{�D���8l���R=��k { ��[�w�w�)�8li
��d{�<ְ,��|��q:®�hK�Oa�:ǹ�#z�!���i:��k/�3��+���gk��6Q�n`�U�A]��t���s+p�*{�8���F�S_��2��>H�Q�(�=��1�1��p��0ꕁ��J�Ӹ��8��hX��İ�?f8�/��%����F;e���͵��z �T�*+��Z�	I;��8#T�9�����K���ߖ�V���<�[����+)��J�B�v��GQG�t��^U"�
%5$=�>� �v5�b�M��z g�#�������a{�=�CK��N����*�K?�B|�ڌ���C@K�P�^�z��4"�N��:�f����1d��/���?�fy^דq�B=����n{<Z�Pp�}i��	��t�I�eY��;�Y\�]���2z��\}���1�L�5�.�\� �h�Jw�qhGU��]�1̇fF���|L͈x�3������e�,����2Z�����{A����C<J�%��d/�s<�lQV)z�L.����Fͺ�����_J��b��a[�A�6H�.� ��9�Y3>ׂ\�Co�����b�wC��zε�q�Q�B;�]{ۃ����z��=�X~�(
��C[n����v�'����V(����Vȋ9m�;��9����B&�8�����\�c�p���5G�jE�z?5�'�6R�Ԩ�)B_�zţ�ҽhGA�[�N��+#,��5Č�s�|�7k�\�|W�R�{4�<�����q���灠�M�[y\~���@=6����E��9�qd.R::�F��KB/g��\b7]��5=,�/3�?,Ŭr:f���)E�a�nY á��(l~����>P8
>-Ȳ�\L�_�)��ՠS��:��(�k��������VF��������0G�@�u�W�`a�ǡ�����UX�,Cޅ����Q�%��*�3IՔ�-�K�ПtA��w�۬G]��뵤��@�K����3��s�R��\�6}��$�՞W|��x����g+ĸ��8v>Z�x�ݥ���c���^���,��!��SkL��"?A����G߸2ހ��V�Hp�_S��������L͹��yk2lc2�L��y�jM�Z������XOq�]�`U����;E��8Rʀ�8e'1O�w����r�G4�9�ѫ��,E����n�W#�8�u��Q��#y��<��1ٕ��v��n��.l����c62�1^�:9����=@!
=���8E�HyH=U�^��o`6^�� W{ �#���0Oc���Q;��;�lՂ�������� o���8���K�;8�v�mĶ���h;@���?���j��l�i="������1W�/�
�f_��P�%<�x��áU�ukXD��q��	�ow��S��;�������M��xǴLi:�k�̘�if�y�G̏��0ۙ�4ۛ]��C7�	}��'?��`�O�C�v]��s��-g�͢^�����;2[M{O�F<�s٢݉�W��9�^�QP���)=ꎃ�9�U�G�Y��� {(�ֲj�D�n�C��
_͞����;<k����9�OC5����A7�1y�)��j�M�C�/��c�&���������?���8Hn �A��������|q[hah�Z���=�T�)��ӡ����/C�w��=+�C�Bϋ/���� ��c��Z�N+�z�Gԏ��h�F���\#�(4ڑ�ht1��U��K�3�ɗ�AF�Qi3F����c�1͘A���lc�����2V�7TF�l�<	W��6��m�}���!���-ی�=�^mȎ:�{�"��b�,5��
������|�W�٣�p︧���=������=ǩnDz?�u��k9.� e9�Ʒ��5p���َ��H���_S/���( �N>�К����o�!c9n,��ζ��#.���g|��@�k��"���2M3��lt���:h�t�浀%�c\̗�k k7�;�@�u;�7벀:/N�,?B�W��w�<W� {q�yw�О�R��EJ-�,�F�h`��g�Fg�w&����>�"�D�E��}���g�Ż����V?�?�Oc��-�;|;�	{��p
�g�/cG�?BC�5��^`��C�Z�l��^�ob/����-������^���{��`/�A�l}��[�x/��I�lu���gy/��Y�BD��?(��
�S�3ɇ�+�G��Ƙ��Xn,?Vk����+������c��a���ѱ��	�ɸ7-6#6;6��ؒ��تؚ��X]lKl[lglOl�P�h�x�ɷ������~���	aW��_��A��_��~�?ܯ�k�OD��8�g�s���"���w�����oB|����m`yHo�� 6�?��y��I��C�xI�����'2D��zɈfd3NF���_�KFی�3�1���g�$^u�;6(�C���,�'�2�f���18cHl�'c(�t�1"c��1�ʠ�2�gL�Y'r�fL͘�yX_���Y:����m����c��2V2]���9|.6�ya�X����z��z	B�u�#���3j�ن�~3v��g��89��ᑌ���L33������\���0�C\�U��+���K33�ev���z�l:D}$]s�`��6;�z���]��)����gv�����)Y�����~P��ř%�TZj��Y�Y�9,sd��̱�}�.�fN>���x��>�0sZ�u����:]�9#q�9[�}�P�%Uי���s��<l|�<�z�\3�޸�M��K�v�{�0U�A9�v��$�%s9��{v[*Va`��u<L���U~E�����$���x�m��Ƌ�f��&s��<���ߛ�FR�S�k�~���A}J�m�^mm��/�:s[��u��9EX��&S�C�#;c;��m*�eІ3�Ď��q;�}���i��c�7lK�3K��C�G;�<��;�0�ߩ�β�"� ���̬���O|fd�	�^P�<�p��>�Sr��5�GVQV��~Y��?�3�n�ʲ*0���/�*k8�+�:�e ����d�˚�5%��̬9Y�e-�Z��:kmֆ�MY[��g��ڛu �0_���o��$�jY�2���>��N�c�Nd�A�Կg�A�l';����*>���-����ǐT[NSǿ���m�;dw�jv��ٽ��f���������'N��=�}|.����,{h���Q�cX��=>{R|���N͞δ�ge�m6���$���ًa+t��,{%�x0�c��^�|eo�ޜ]���)>{w�>���GأM�-?f7d7���`����sr��B
s�s
Y'9�r:B7����:��ӝee�rz���@�A9�ɺʩ��32gt�؜	9�s���ș�3/gaΒ��9�r��ϩ�ْ��e�ٙ�'�����?�P�ќ�9M�6�_n$737/��=�	A�<��
�u���6���u�u�RωYG\&���Qzn�ܮ�=r�r����oNg������0uޝ4�f]��a�����mF�K|�����!|�/�uA06�9SnEn�
��`,��[�zȭ��;1w
���v��C��������,�j��!Z���$�������\ʫ��
�oٛ�l�M|�ϯ��[��q�5�˯!��?�xG�;�v�܎�=���q���f#ǭ�8n݆�+�w%��A�;w:p�� :O��S����"��o!�Ŀ��Rė"����H߈�w��{5ҟD����E|.��#~?�W"~%�#���� �һA�i�w�k�^�qcǍm��8ׁ�cA?�jȾyː��{���3�?�@�/ ��{8�i@��Z���g7����<C�.�u����x��V ��[����A�FυA�-�ۂ�.ೋ�/ܽ��ϳ���>�&s�.N	Pֈ���g)��o�·����Q��H�٧+����� �7��*(�
�B�/D�T�OU���5(��H�5��>dD�1�v��!eo�˱P�rM@�	��<�=���Hߩ�%v,SP��H�`G�;�qnC�JH�;�r/Rf ��I�
��WQ�WQ"ښ���|�~��#�z��u�8�s �7!�&H�]��.�#~9�|t���yH��8ڋD{����?#�g���dn�o"�pz�A�И���"�,x{�=:�����`-���C�<4s�*8���|,8�8�m�[�Ay4�ȃy�Y�ň�A��ՈW�ׁ�B�Y�Z���m�D{�{��Q��#�>�O�n�nDY��%zxs,s�Q;����/ �|�ц�p,��UH�B��V��A�����R�K��Lh>|6��&�â\X��EIX�]��H�!/zW���UHX�=
��P.zN=���f��Y�,�P·@�CH���!�3�;��(x��έ�s+��� �7�{����8�я���$�/�k9�.G���^J��0��"�/B��{�	�im�+�)�f�v�cEW����&���F�D��xYԋk�6r�3�i����Q�'<�b�f���牅b�X.VQ�F�'�Jԉ-_EyW��������E�a#��3
(��hot2�=(^D����(5ʌ
��nT5�8����D�)p�+��8ya�|S>����HK wތ=���`hahN����3��q��8�:����^�7�^�C>����qs��#�؟"=���@����|^�k�)�ĩ�C�w���0�y8G��c�G|2��N���]�3�)V_���y��=��&��x���<����ⶢ�h/:������K�o�Ţ�c��'��/�[D��M��Ō�ߙ'���+��:�G��N�
Q%��/Մ9NLSD-��x�6G,K	���!���%�#�%2�{�Z��ҩ<�4�	�����G ���!E��V{c�.r~+���b�΀�@S�^������hkt������o<�����p�کq�9�)N�3әCn���Y� 8�Y�u68����;�����v�9'\�Lqg��t��mM�n��u���(�����K�ǁT�pw0��T�&;w�+��**�9'�s��#(}��aZ�Nr�?É*�����"8E��M%	�o�b�;�8�O|�rj��9T�\���	���]�.&}� �e�Jg"I��m��?{��YK�׺�1uw����D2o���4��f����t�0��3����$��܃�S4�����l��t�1dr١P�G��!���&��;���,m������s������P�f�7�t�x&[����0ɧK�JB�'{N�ZV>T�$����C#����áєlh�;����L~ZhFh6��B�BKB�C�Bk(�z��)�=�<ه�(ߖ�6�uN>�3�ǩu!�?t(t4�0t�YJ�xm�����3[�=�� k	�PTk�6���� N�����.
�	��������^6�=	�:^��ܾ�#X]�&<.<1<��F��?��a�o��9�I���9d����Ë������NmxCx�7��a���vgEx��(�7| |؝>�ZQ�DD0�n��5��H4�i�l��v;D�F:D:G�EzFzG�F�G�v樖�z授��K�!
죑�n����"#"���jkZI��-F-E�D�s�F&Q궍LEn�$=E�;5�Y����őe��2�\dI��9�H�щl��GvDv�}�'EF�S#G"�F�ty!�w�z�^�W�#�ѝ�uq�^w��W�x"�� �ܫ�24�9�/�F����Xo�7���M#Z3���<
zK";��|�[��V9��z���B=�Do�����}���;����{M�M�r��c��MQ;	���Y��ПR_LZp��Ѽhi���!�&�>���J�=�]�E�>���[���ҝ�hE�
nx�:Z����Τ6�5:G�A6�5��w�>�!���Zg+I:9�"ʧ�>�@s�;�hϐOæ�
��w!}�>¨>�|�Ob(s��61��)��0{3����L�fc�
�)c�
�řnu�앯��j���:>���k`�.�=��EJ�kF�������9�r���~��)����,�Q�?{��ڃ�7��@�*����d�֨�U_;���b ����RpX��+�qz�|���QE)}�Ƭ�|��1L�%h;�b��1(��C�M3'ޙ7)�SK�,�z�1P���ao��&����Rv"e����Է���N��[�9;��f)��;��P�g(�!]!�~)���j`F��<���'�n5��~z@����k��M��c�����p���?��k���;(;��.��P�	k<,��4?m�k�[��{σM�DY�Ҋ�SN�n�U������f �t�j��,�%�-�f���I�Xu0[�r���0T��Ō[������bC�oy��RlH�4:%�}���0�;!e=J<���p�5`>�vCWj�P���`WE��U{�U�����(`�w�Bc+U���-@JOhi8�e#�����9e��N��؍m��(�,S+��G��iN@����:�|Z��W 6!��fV3t�KN���i�<���s�	�� һ��e�8\~����N3�p}uWO�U���h5LA�����_�~�铘��
p(�o�ɜ'�w8�`c�ѷ0�&��'6�N��]�?�n[�1�UX��	�hO�0S�����[륮�hd��Ft7v�у���t� �#��7F��L�!�>�\���ɷ#�Q��B��{�/&_B~ �A���W�F~$���ǒ����������#�PǗ�����*�kȯ������F������%�u��!����I��S|�K����w�ߣ�ܯq%�B�Q��5����Ƥ�Q�=�wI��<����ۺ�h}�.��*u@e��Z�!�]�<�/�C�y���I!ه_���ɉ�1[�~��e�H
�h������%�~)�;ig$�Z���]�� _��g�,���y��#}U�߇|?��٧	�}���:]���Sɟ��$���4r��ܾ��,)-5p*�W�N�:M�^��z?۰��Suw�a\�3��:�t�0�o�0��.)���~��E�m��>Sx���~���;?c�Z����I}@ڐǎ%i��6r�6�v��aj�r���LaR_�6<S�AZ?A��>y�ܒ��������:�7Z��ݯIؑ?.��x�N}�?1���c��D�>���Fu��c�3�׍?��|�t��	�K�jJџ�B��_�\V��P-���&�[�o'���^��&L]�E����G[�����S���5�!�矈��	}��<c��j�)��ᐏF�m3#�|+�:��!�9,a'm���ł����et �Y���E�4�=�������	�2�j[���Q�Ɨ$p3*�2��y\��g�~��h��4?f�����cȏ�&���$������%�x�S�t%+˗1��\�As]e,&���J�ϑ_G~#������ �[ɘ�/����Am.��aF�����LS�`Ίr��,������:���˱Izڭ��M�g�}dR]d�'��X��S3zc�-����m�u&��-���$������y��������x;�s��v�V`��V3;*=dR�dr��]�Vr�/��*�V���)'�`h��XOaho�>C�W�[ʯ!� `G��xC���u�D��N�<��{���R��<��W#�$�\����� ��NC����)��8�q��{�>�_��#Hi ��]�?`)�o�)mA�(�B�d@��q�uМ���
�Bħ�)�=�!�l!}p�G|'�_E�t>����=R ~0�x9p���<@�����o:ȋR�gA��@�$r�@�ͱ��[�A9)�� V#}p"E�2tk�A�G	8�ވ\�@sҕ��#�-��U���A�_X
�3A�	q�GB?v9��.,GB�(䅝�м�v>��}�w�(pnE�w��#��#����� �a�/b(����c�0E�Y�n�3o����}�����g�gć�W�"�����nw���=)�O�F^��(���G�EWo�7M\���%�E��-�G�D��D�������"!�I�
���0f��K~����k�+�?�t�~��a���f�9���A~�N��㌻O��?B�A����7��LŇ���L�Q-��Z�g5�w�"�Aat6�=��F_�����?c7������r���1g<9'NfO�3��,c.��bc���4�ϱ�`'X^�s)Չ���f�jæ��cO%����rՎp����NY�,�����}��w2?����t��8C�8f��H�=��ن�OI�é���M�MD�.ɇ�I��(���ܗ�z��}�}��͟�?����ܽ�0�%�h�M���}�h]]/>�� :\4��&���E��ɷJ���im�w �9ͽni���{��M���x��1\�OUU��P��ۦ �j'�$����J-P��أjN�;;��(��]eWQ[���S�j�����������õ��w�]�]��}�}���}��u��~�~X\eϱ�n��Z\-�U�	w	Z]��U�a{]�'�uh�&�Y�6a�;��U�`�����4nI�<�[r�nU�&�[��եq[R�6r;S�r�ӸC)�(�T~��K����I�\$��L��������@�q-]ڼmҸ����*{�"r}(�i�ҸRY&+d�N��b�]�8���&k��8r)6�\m73�����O�Rq�E��ע̥ri:��+�;�]�Ɲ-���:H'��i�Z��<oM㶧q�R�^rR�ar�R�[�F�'Z�t���L��G�d&`w��x�{;'Nb/ESq��<��j'@���{PԾ[a��q�e�WT� W�w�������حbm�V�kw�wՉ���4��5��E�;Qo��N���}?p��7�z�	���o��>�V�*D�yԎ��&�e��|��=��zN��a~U�6Z����~���/�O�����?�i�#0:�!�K���Ǌ�N�1:= $��-S1Z��9i���Y�Q%L�y��$���H�"��D���C����^�N)�V��:��>�bU���n�1ǘO�"�K��j
�S�����M�V\o'���V�{�p��cO�LA��?�����v�m�t���u&ߍ�����I��������쟐��H��͞"��e����������9m�"��`��ɽ
S�_88#�k$rqz}��n�?��t ���}t|;��#eR��8�>��� [�����v���p9�\�g���8a���|�ZG�b��Z��-r�z�G`����՝D�!�`��(�y�A6�U{϶�1�p
�yG�%�\�o�3�O�t2�@Wу�a�z<�����is����1�s�����W�}����UB��D�v�#I؝|/Q,J�&J(m��x����#Vr�5m�Ω>'y=5q�G��0:�Ғ�6ћ������(�'3a��*"ޣޣ�JiVi�7���=on��Ϳ���_�%��L��$�7����͂רh)��|m�xN��<��bN�n�vS��Kn���-�n�v�S�sک���t�����l֛;�����nA��e���%4������i��|�Q9�W.���Vnsׂ�@��wV�9�/p:�*Tz��Zo�����fz1(�N�^��O�wzsg�d�5��N��p]�������N�[�p%� ��enB/��`�m�I�] �t;����5�K��M�ۄ1�	s�w1⫹�걚0�6uH����2ܟh�j���DO]JF|���fOR���
���-��F��r�Hݬ�s+��3Q����#3"�E�E~��IdA�Io�7K�ȥ�V������T��Gk�ii}t���Y���q�K�-��n�X�� ���5��2o9��I�k����-�*|��
��q�-p���%Q[��-O��SS�|�K�\��`jڮ�Yn��=���bv����e5��;��5�{��c8_��+xl}�!���|�|\��3�l�YaQ},6��L�ƛE5�q�:��h��f	�y�\P��h�kWzA�EKQṞ�&��cB�"�4�l���P�'�g�z�����ɴO�A�E䠾�M%����;�?�8x�%��ʵ=T�e\�r*he�f�U��\��T�pQlF��R�e�z+|�z���50����H?g�^x��C+v�ȗ_�.���_T˩���S�-��"[N�E���4���R~1��������.��|�7�,��2b�$>������'i͹W\A뤿���ᕢ���0��Y���e�DT2��F~�y$������Ȝȏ"?�,��,��$kj��T�yH���8���.��Q�Etyq�O=�-M5��}_�9��r�O���'�/�x׼-��vn-b�h�Vn`�e��ϭ�<
�S�ަ�ւ1��d�����h�q�����h����L���uY�����Z���(~�M3�3�K�砞gby�pͣ߰����=�OZ���ѳ�䇞W���p�tA��{I�.H+<����4����s/{�^������ǵZ+Vb�X~�j�\y(�hM��|F�������g
��<hH�S�5�s���.N-Կ�P�����A=��/�g�O~��K��(��$��|���&�{�(>N4���݅�����2��;7�1�1q3���e"�$�S��C����)4��[Iq'%o���;�n���A�Gd�ltL'$��q���u�骐`;��.��wvG�^�S,w��by8�r#�/���� �*�=�DΠ��8�h������P��a�SI�S
]����SRg�3�p6:�	g�ܜ��F��)d�	6P�X���J;B�8�ɲ���Cj%��#��a�i�'WQf��A�4E�#8Cq���]���ɧ�����9]�����T�	���ہ�v�g�5��o���g���ʝ�"��r6��#׃g�G%�ՠ��;���5�lq����G햚OSu�yg?k�9�%9[�p-����I��N��µY.7ByV��n�$M��td���g��\{���9�n��mﶡ�;]<�mi�gc�ge���:�dnW��[��q{����/�pˈNG��VF)��)��
©b��Cg�[�:���n�.�1�zY.����h$���D��w���Q�%n-�Z����O$��S �������K`��`KTD���f��l��\cYÄ�Ι����2�Y�΁��p/��R})Y�>��U�.�;�Fܥr�����]���]K����t]�S�֌�I�Y���A�n��G�+{�Y[�����=>���v��ݻ�ѣ��S���P�q����L�P;}��^��G�P�)�n�OG�Rg����h�����.f����aϯX��Ԟbuz�ډ�v	��.�:��d|��A���'R�R-����@�䭃�AWu���O�B)8+���xjo%���Wj�O@�:�[����ۭ�a��l;��=��N�V�`'����Y�?%d7��j�~�bP+�W7=��9e*�Xx/�O�����"x�qn�},��,�<��dEB�^T�J�dJ�N����^����1�[��T~�$-r��M�������� u:�,I~\u���ޑ8�R[Rޒ�^`����[E�o]$i��������B=�j��r�g��~����?'k����������\��ޓ�II�"Z��g��O�JϷ�����L�@j �);�=���J�@���I������g^LZ��s���U;y��i����|�N�8�?~�:.G�z��:~��+��} 8
F���k����Q����|�S���(��/�~�7V$i�����ʑ�E�[\C�~ xr��T�=e����W&l�۱�gw%�޿���E6��?�0��4ʛ�Io<�M����(�JL�\�ϛ�b�2����K����c���X�		y�0�߲��U��7P�bҿeMr=�[�M�ɩ�-��w���*i�kYe�zy�����M��������ƞg�[��֢��X^S��̵�b��m%�}�s��۳�';�΢� �����Ss�ty��1����l�����q�w�]=��y7/)��|`տ!��`�ॡ��VҾ�KC���U��^������KC�CHۣ	w4?�h���66�'�¼$e�ڊ���օTB�E���]�2p[������cw�/��B1*���ґ�����3��Χ?9۝�������9N�����tO�.���������x�Yn�)`�}�upl^�O_�n�,�Ad�~q5����^�x�u$��g`4)� ����}P�]�%���/�vWɵ��K�ݝ�����Q9Z�3ąz�t�G����q�/�\=�*��ִ~�y��n�sGq>V��|��Ns��ke�j�Oӕ�����^��L�&�gI糛��(�mO��.Ğ��/;��1Y�;;�MG�����]<����h���c�Ĺ�4��a�x?v<��V�7�����o��,6��q	p�|���.-'s�~�8='�ϟ)����g�5��Q�|<���Iг��Y���|ڽ1!x:�|���AQjTU��B1� �k����"����ٯ&��R��^?�Wfl�p�^QF��9�2��V�}@S�]�y7ٟ�?����׼<����1����*�y�Dy���v��E�{Ak�q�(ϡ���x!ZBݩ�����O@W_J��7�W��H��f����J�]���R��J�O��߁�o?��^��Jq�����X�$���k��������7A���k^�೐�9���9��E��Z��-�f��s��X���2}�8��Ni�l����C��/���[I���)��c�x���EcȬap�X@��N�+�sb]���։��-���y�U�����:Tߧ�Z�[���V���+a;��V$���k���K.����#A-�ӟ4�(陿ʭ�7����EM���8�2�S�oe?�����~A��p�Z�ս�b��@)���J.��H��n�3�����A�*�σ�9�h�� �]E�2@���	�i��V_�������������	��h<��i���;�7N��E/�[%�/N��U"��w���=���P_?|�������JG�ygH<���g�8�/mU9�|�,�L�= �g�W��W��������Y������I�Ϝ�J��nY�-(��=r�r��rO?�;$�}�i-:����E0���>�����B�Y�,����^v��N�k�p?��G'՟t!��u*�_��u/S����.N�6��&�a5Z�^H���~W�S�*.�7X� �����AxV~�J�=�ex�����e�g�>i}�E(��Q���
���9��P��#�o��QӘOZ"���{�GC��r��X��(��nK�G�YCZ���������4e��s>�Ԝ��?�����9�i�m�S����8_N�qk����R������r}%ϩ8C��sg�Sq*���}��Z�ܕV�y�S�����RӅ�4q�cݝB�?�bM�����i���`���CsoZ��ij��5<�-������X#�p��ki���sſ���i�W�X(j
�4ܷĪN�}K��H�}K�Qi�7p�u+�תo���*Z�Nk-��2Z�դ��Vӌ�}3m������[�ݟ��[�M[����ߋ���f[�K[�-�H[�-�Ƨ�/����Tv��4��Û���tx��/���"$̓�z�~M�Xh�*Z�'_?��������.'��yL}+�#d�� ��_��Z�#<곒<_)���-���	S������ct��lM�-��UC����mv6��I��ٛ\+`(���o����`��C8�q�b=͡�5�RFQ\�!n��Rl<��x�f0Q�$U�
2?S����=����i��Z�d��-$R4��҆�m:垥u��R�-��n�y��G�*e����2��E0K�S����E0oӧȩ����"������d4��I?���p�����H���?��E�����8]z��'����v�c`���������K�u�IՓM��T=�RO�В�ڒV���k������9��-U㜅��D�,��]9���6�_�+�� T��a���<H� �3�#k ��d|��շr�|�UHX�e���3w������^�:���GyJ��,�;�̲Y�f�UI�J����Y�K�J
��as>�0�S��0�9�:=N�T����tzK�ߝ����r�z�~��%�Ey��<��[#�Mt�Z���L�Iד�i�2���⟳3���to�5���#�%�ejB.ŗ5/h��D��Aߚh7�%�6��V��?������ۊ&���9��H~���x��wN�׊D����f1`MR?�g�&�f��9��ߎ>C�i�?�Zx"l�4�oy�C���*�o��O�t�m@=���Þ��a]u�D��?Fm�Is�������4���W�?�;�ϡ�6"F����Jo�o�ٷ�󤞵����h�'���b<-N�<�Z���&�ӼN��<{_A�\��A�|h����H7���o��p¬:CV�H{��>s�N��e��7��\�s���0�_%�Yg�&�[�8�*���o�g�-s5�U����[�qZA�߹�������Ex��	��6��Xq
�J�<���e���Xkl��dlE9��Dc;a�+������q�^�@0�gԝ~��&i��.iܚ�:��e�K�=�|Mb<Sg�s�ՙa]t)'S���>#X����g��	}�/q���g�j��"z��)���L�������-�b�`������b���A�(|*�$m�Л�.y��Ҥ��wL�h=�\n6�D��x�F��z�XH)uz�ق�mt�c �ϼ���zZC�;�c��ޞf��c4Y�De�8D�(譡�㢉��Ae�a#�Ȍ���'���GYN�?�wIҤ:q{��U�lk�|���L�Fm���i6>���s�ڧ�OEq�'xի��$.g��;�~�Mw�=K��+C����ꛏ��qգ�<Z�����D��o8t��'��g�>a��1c�[^0��C�F[ْ��<�*vu�O�]�vW�D���h�Ɣ�N�J��{-�\F{��ѕ�{,2�(*F^�}�N�|��Sٷ%�ie�X��U�Q�Л��,̯�jުN�6fSz�X��ъ�n�quһ��۝��v-���^^|	���݀��?�4p>�T/ �-��?���4 ����ij\/����� �G�o���zQ���Ȫ����-B��k���(�}�O��I�#{KR[��;먦���j��ڏgo`���vD��^�[mޛ��VW�:�~N>Q��֠^�V� m��������`uǎ1�X���5���ǩ�Ԗ�\�ڢKZ��[�@�rms���mMeK�Yar��ejnx,Q�ɳ?��wQ��NҎM��2�S5��\��=Dbo��jI���QQ(ڥq���z6q�J�Z�����+K�E�3�'�R,g����윟�� ���s�����j�`�����N�H���X%�:�ɸ{�K��?����2n�
�����z�J�CW���� ��	���*a�z�O�ecz��Y��ax��{����9�an�V6u-�D=�����o0DD�#�ml�1*�w�7��2��rQ�&uJ�Է��Km(m�FS�EI!���F��8{gj������6�,�`�ܴ��K�ǒt�G��]Io�J���y�R��,]����L"E��i4U�V�ʚV���V���������qaZ{[�V��RRZqİ��¾sԝ�"�ݕ�ĺw�)��v�����u�������T(Jo�_\(F�VJ�zѓ'�~�����4vW���'g94�����S�4�]��Q�(2�eD�c4B�y�W�x��Y��,�J\N+�O�O�+D7q��g�0�����iV�{��=�o��[�O����+��ͅ�/�RM�Ģ�3qlZË^w�9b�Q8p"��ڻ��Z�1p>�R�Հ �24`0�jĽ����v���`������,,� �~��{G�Հ5�� 'N�����0kg������i.|�p;���5�<
x���eF�vwսV&```����1����``�QT������
+��.=��:�T��{��ݴ&[,$�jCVҖl��Q{��dM�:�-v&��VjG���/�x�;�>|�!�^X���ϩa�i�(ɺs�����ze���m�GT�T�_�]��^vZX@���4�]#6�]4�k4�4o�h�1fK�5�fc�q�h4�f����i�3��V;��l��Z�����2S�βH�Cd�� ����,g��ʝ��t�Z�ڇ�����B�BcBSB�C�C�Cu�����P�U�}�{�o�,<,<&<%<;�X�����ùdS�5�%<�����vI��c����ڤkB̜�t��s�z	z���)�شK�V@6ܑ�Ξ�yNy�V�p�
��u�W�5:\��C�mRј9�:����H�j�O�*�^�r�zM���:5������9�\���|�6�~Q���)׊^6��.4��%�T���p1J�i��!�4�]�$n�Z�[uؠnPa����*���n��p�
?>A�U�	S��*l7G���Wa�v:\��O-J���:l���J�k�ð��j\�ԋ��s+8�hj{�9�tؗ�J���o���j1FLS�t1[��im�Z��U�V��Va�q�
�Z������~MO�ԧ������g��?����S��U�Y�C����*�5�y����^��C��h�u��ã*��H��txH�]ǩ�*]�W����h���\�WM��r=+�z]�5ѿ����kV�\�5�����_�k~}S��m��^�nE�^���o߇���F��E��%�Eb��׊���.v����������P��~STxs���P[]m-���p�
��k���v��R��T8��a�ש�M��o٫�R�{�V�p��7���E͵tk�si�pvzQTt_|k�
j��סn��ѡ�u��b��^�Z�2���t�C�_�Cm냵4����Q�C�K{���Җ;����:�p�DN��<�mu�5�e-S��B��W�,_�e���N-Ý�UXY�|l�L�)Ry0i���#��]���cIe�XB�*H���\檔���s�uY�����vu����#ͯ��N�^؜��[��3tG�v:to����~`����C)�k~}�Д�CI����l���"��9�K��2K���3o��-�[�r�p.l���!�w��sw�;E����#._�#
�υ7���"/�+"��z�՛�MWE+�w�nѻ�w���5���5��F+>/x*qVg��3L^͆��V��hct0�=��F�Qj6*��b�1��bL7f�E�2c����H��m4��Gs�c�s�Qgl5v{�Ǣ�h2�7���f;��ٍ��$�@��V���Q�Xs�9՜!
�
s�9Ҭ1Ǜ��i�Ls���\�����Mf����k4��'��5�jeZ�Δ�Ѳ���kXm�V����*�J�2k�5̪��X��V�5˚g-��Z+�5�k�(��X�%�
�9k�Ugm�vX{����j�۷���v[�����i���R{�]i���E�z+b <1������n�H�oE��#.·#!�'"4����:N�·"Q��#1�oG|�'"�}<�IWov·"��Gr��Ex"�!�~;�GW'�2�oEZ!<�0·#�OD>B�'"�!r������Z�B-���!�FK�q-][-�'�t�\��r��r}J��A��i��Q��-W'-�g�\��\W@�.Z�+�\]�\Wi��i���\ݵ\�h�zh���r��r}r��r}^�^���:-_o-����b-�Z�>Z�/h��j�n�r�h�n�r��r���k������E�U��r�rݦ���]�U������C�U������B���5D�u���R��]Z�*-�ݨ��Z�{��ô��j���õt_�ҍ��}MK7RKW���-�(-�׵\��\߀\5Z�oj��h���r��r}r��r=�������k���A�5Q��-�$-�wu�M��=�ڛ�����o���a%����Z{��^,���/��ЇV�iN0���4D��lZQ-�y�:�Il���q��쥵~o�1r��F{�{}���4B�u�����ֱ���9�=�c7G'Rl�c7G'!�x�ձ������ӛ���8��qz��M���~��,��w�R�c:vst6b�(�q�9Z/��r���}$^�x�?��;3^��r���}"^��x�?
�������k�Ⱦ�k���=��"}a۟��3v'��o��G�F���6�=���[�I?�F�m�ʮ¾�N�5�Bڏڏ�����g;��v^���3�+����Vy�<N^�_!��~��>4�2,&v���*��!�w��b4���/��҂Si��6�V6�3D�7X_@���;�e݈��p���qwp��1Px36�R^�?A�h�K�P0�q)�y;�p)
�<��L�h�O�-���1��/[4�F�(��^$�Ǿ:y�w��~�=����I�'����yg$�ΐ{�9��ڕ\G����\r�-�һ�+���F�/���%����s݃��q}*6�Vر��z�T�k��)����fùg�o�}�דN�r^s���>G��xJd�_�yjZ����ǧ	��!���R��Y�Z?Do��~��)Lc��m]M��<�����jG��O�Y�I4#�bM�Y�tk&�L���t�N���t���椫hV����M����n�v[{���A�u�f�G�������+��]�n��������}RҒR�ғ2G^&?"?*?.?)?-?+��W�k��s���:y��A~A�(o�7�/�[��vy����K�#�_��!�!��o��$�=�}��|T>.$"��O�_�g�����o�o������%��|E�A�Q�*�$�"_�����1�P���@o�W���{�{��������k￼���~���{�{�{����'�/���_�7������㝌ZQ7�z���񱉱ɱ)�i����������ؼ��؂��������؆X]lslkl[lG�!v"�䛾�G|�����|��o���/�/����_�ؔ�%늬�����\�糮��B�Y����>n}�jg}�����
�*�A�;�w����Y߷~`��z�z�����I�)���/���g�g�_[�e=o���{�E�e�֫֟�׬�!;y�����ֻ֛�f{�]oo��d��>f�O؍v�Ҕ�tdD�2[��|�Z���d�Iv��dw�C���d��-�e�W��~�� K� 9XV�J9T�#d�-��qr��@�7EN���L9[Ε��B�X.���J�Z��k�z�A��Mr��"��z�Mn�;�N�[�{���]�p��
�V�6�K�|o���[�-�Vz��5�:o��ѫ�6y[�zo��������{���Q��;�5EͨE#��c��}7�P����c?��0�X�؏b?��$����b?�=�m�w�b/�^��1���۱w}×~؏�Y�����/��o�����vG��3^���5�{VϬ^Y���d�d�OXmhm�Z��ag��u̚fͰf[s���Bk1�W�zp��ʹ�F��]��G+�C�\���u��A�a�Y�C���r�1�	�)�y��J�&�$�,�w�޿*�_�ߔ�"Z��;�!������|L>!,*&.�������i�$������]2f}L6:±����O��y?���~����O�7�o����?x�z�^������w�M���޻Q#*��ظ؄ؤ��،ج��E�%�e����M�-��������X�/|��Q?���[�����?dl�ؚue��Y�f]�uC֍Y���$�Wv�=���������ɾ�Qox�4�|��3a�d�����X�C���Ƕ�dw	��.�>f]feY��)�֕�b�a��1�	���O��Y��~e������%��֟��X�[%ͽA9�ao��j��(<,C2*3e�l%d�l+�ˎ���*�2Y.��*��p9R��5r,ѺLN���TY+g�Yr��'�Er�\&W�U�9{�\Gֶ��.J�;�c�Z�vo���[�-�Vx��缵�zo�������vy{�}��w�;���"jG��ož�N�{�Gb���={*���3����>�b���b��ފ�;�[��{~���_�����o�x!㥬.Yݲzdeg����iq�im4�q���b5S��[����y��1[����������}B�����&��q��	�D�jE[��-J�����)=�8ﰓ�F��xI�ʛu'��pZ#�i�)*}gW�����T�/t�ԗ�z�ȳ�"�͎s���)��i�9�2^bePb�\��B�؆��-�h�4��Ici�4QL�R��!f	~��3ejO?��4��_R���I6NsGQ��ޚ@y�QΈ>�rf�t�b�Pg��.@~S��<�s෨�����0��[C~��O�N��"8�z������մ�z��O�� �w݃O�~)L�#=K��j@���{y�����W��򾁼+�w�u1��w�À�x�M����`��c�~�kb�m��H��z�m��Ԛ�ʦd�ʷ�E���u���/�/�Z�.2������x?$���2��<"
�?�1�F6�㢭W��">���~,>H�ȫbkc���b��I��?������7�7�7�2��S|)�北��Ҭ��S����K _ܧ9o��7�	H=N��^��
_�Ǟ�6j͂�M�Z�����z�QR���{R��F-E��Z-��Sr�VR�^F���m���vR�1u��_.)i��2�`��Uk�g�V�D![����f��b��-� :����#"8��%�ֶG�����	�B��^���4�w�cZ�DΎ,�޸BTS�����)6F��x�����z��<dP]�k�ڏ����Q����Hq��Η@m��AB��r�Ә���ET]DG1�<?cJ5�Q����5*��J���Z�e�8A=e�K'�(�S��1#Wl������]�����e4�I}nO1 3�	�p�"6E�P�X�a��j��ij���Kuu���O��^q�Qv5L��ɱ����㒩�3��tv�K�SI�Ѝf}ݨ.*�8��n4�,Fr��DUCE�����#���}4~t�~�F��M�W�a&���x�Q���l��Z?\���p�z{ͣ���Ɛ�uA��X)�i|*}�j����x�\8>rH�4��.���H���j��C�Qp��x���C��搾y\�J��3�H�}�o��U���5��k��e�un�~��Vۥ�d����Tj�m���_u�\U���s���'���e�d(c'u,����<�Cd|M)C#��#��M�c�:�#�x!!bH�#��h#"U��cċC��9�R�o?�&����ė�����s�9�gw���sv�x���͇�v���&�_m�7�ZJzcj�e����/������m��
���G�s���Ǻ�Z�}�o�E���E;��_}�J#�C�W��#Z�����=?�7���ⳬ���^oM����Gb4�5��j y=��_�(����LV����߇�x��it��O�6��K���S9�1���q�f��j��7�����2�P��/	����r�˫����c�ݓ1�'�*n��sOŰ�f�H�\'�^it@/���S��炃���Xr{U������P�4y=�ˇ��vC�:�3].:��ĳH�k�K3{'%�İc��̔��_�D�wq�|��ryO��U��s������]e/}�W'껞k�z2����G�k��3z�z\uIH���J����^�Q�G�J)/57�R�0���`�%=�KעC/)��=� �3콣��/���\>t/^w&=��1�K�Ԩ�*�x��^��uF���W������Z�l^OA�6�o�`�p~�#�=M�`���NԒ�-�k�V�-�@�̠�	��%� /_s�B�W�G�M̔}t_V������Db?���1�ƨ3��<G^�R|���L��g�]�_W�7Үk��%��Q�/KX��LTb-�c�t�ZT�֢ҿ�>����E���uU�^}A�F�[��нU%9��_�Ub�%gUx�/�H���SB���D�}	�ΗP��-�hF��_�_&=e�GIB�^����|	�_�]�KX�ӑh��Rt�/�C��E�/*�xQ�ɋ���EWk�~�_/Z�7�6�kD�H�]�k�a��C寗r���Q�A�Z���9N�J���1�:�����I����d	md\Bz�N��Vu��2��J$_����ա�ІPShw�9u�R育T��T��P��Ft��T�J�"����ݪY����V�;��w�q�m�0G��)f��k�Ef���\lF�
�ڬK�72���f�y�<o^�,+�ʴu�]�c�ZV�Ub-�[Q�ª��V���jf\K��n���[l�N�3�A�P;�a��'�S�;�.���{��؎�����qi�S[����j��"��C.�P������t�$G�Erd�\��5�cM;ޚd�/Vώ�!v��E��<�В�2k���zLl�Uj���s{F��V�U!v��j�V[��Z�rƛ�6Z[��bwZ{�}b���a�%N�=n���ŶYq�k��o���~'���6lǖ���[��b3�v����fr�o��G�n��ǈm��'��()9M�T{��+v��gK�$);�^ v��o�؅���b�O�O�eb��R;&�Ү�kŮ��b�ۍ�V�M�N{��7�f�����A�����}Rl��f�Ş���ߊ���ξ ��p�t,�wn��d:�p;C�q�9w��v�;�ĎtF;r:c��������t�9�L'O�,���'v�3�)[�,t��y�yZ�SN�Y*�ܩt�ŮpV9b��N�؍N��S�v��Y�^g�sP�{N�s\�1��i{�9���������!�G�r}�t=7��{�;�,v�;�&�67�.�Nw�;Z�]�Xw��	�dw����w���,WZ7ߝ��[���>�.r�������[�V��pW���ָu�z�kݍn��M�v���ݽ�~��������cn���i���v�+��_����~���Y��)��2Ħ{�z���yC�fy�y�bo���F����;ƛ�M;ɻ��;͛�����{s�zE^���c�"����Sb{�x�b˼
o�ؘW�Չ���z�n�6y��n�v{{����y�=����=��N�=�{_��{_{��~�}��(�BX���D'��s
o	�����Ya=�oh�����wGxDXϟ�s�Ƈ'����)�ia=�lz87����z~׼�����U.?��W?J+{��V��H�Ry�,�YH9�Ry��9�R�R�R���!�C* �
�2�2�2H%�R	�ա�?��u{/$�A�C�C�C� U�*�*�*�*�K�� /Aj!��Z�j�j�jH�R���C�!�Hdddd-d-d-dddd=d=d=�e�ː�!   �@^�����y�*�UH#��y��5�&�&�&�f�f�fH�	�����
�
�
����������	�	�	������y�:�uț�7!oB�B�B�Bނ�y�i�4Cކ�y������;�������w!�Bޅ����y�>� � � ����0�0�0��� -�H�Cȇ�!G G G G!G!G!� � � A>�|999��1�c�	�	�	�'�O �@Z!��Vȧ�O!�BNBNBNBNANANANCNCNC>�|��i��A>�|��i��C��|�rrr�%�K�ָ���Q��,׽?�U�E�a��0�s5����8���O͏��E}j~4N�(�S�q�HQ����_����h��Sԧ�G����>5?�O����8���O͏��kE}j~4N�+�S�q�`Q��������h��YT����� ��g�jRY	Y	Y	���@j ��Oʣq�xQ�6��ߋ��)h��_ԧMA���>m
�O�iS�8�èO����+F}�4N�1�Ӧ�q��Q�6�ӟ���)h��eԧMA�>m�O�����^��,O˅�Br!@�< ���y� �AH$����ɇ�C�!��4�O���Q~�x�'���uoُjUgѸ^�C�ݐ�!c c c �@��Ѫ=9ec�q3�'��[<ݘ��_����a�
^Z���]<��}o���^�]�y֣Z��?=jI������d=/R?���'(�3	_��QÍ��R�
Y�eT~�QaČjcO�6���Gz���]+w �^�HW�r�Q�����*��~��W�-bfu1+�.dM����?������G%D�2�6�~�K<y�=m�\*�G�������K����m`�ڷ��/F�W�����*Z��\E[�}�Ѧ�h�b�]1ګ5w-U��)F������hmb��U�31ږ�I�6$&���V��ީ��F<t�Jy���Ӽz�C}Ɠ<=�#X=v0�)+��X�]Cw
+�;Ы��l����|�O<��i��Q������=��0�s�k��3oƕ� i�PnL���D��OM��&<Q<1y:e�U�5?$�R��?����^��RcJbʴ>�
�9:֔��cqn�&��xϬ�Rk5��;��=���w>�V��9]x�FR����g	�o��_ح�~�ak��r�vl��z?����U8����rG��y-����\���V��<�ԔLMq���7�}Kb����xGڽ�_)V�JKg�ё9��h�s6�N������q�NgLGo�Q��r}�oP�M�^HƥgƔ\ҵb��g�Ѻ��!������%�����V#xK��nl}�n�gDKx.�)��+n�|+L���l\~��N�$�G���_}<p�h?U�V'�rۢ����:�X���mg��V{��?���U�իrG�W������y>�8ϼ^8�k���١�y�L��n���g�<��<�{4?��l~��r~����\ף�������^�ϣ}�<{�<��y����<�Gγ�G�φ>{}~���?�����{+���gPe�W	=�^2� z��}z���o�<=�����3^�K|�yd������j_��3��f���
'g���>�J#9�o����ν{�NW=r���ū���+H��>�^}4�����J�W�Qb���x�Գ��k���WY�W�uū㽐~���{����sU�U3� ��_���>����:�9�{�)g����R��eĵ�c5�����F��
����w#������Hz^Vb�H~�7��ȜHa����Ñy�G"E�G#�#��,0��'V��s�D<��HyW�(���
�l#��䣿A�9h!�:}��>������ߢ���}����A/�������U����PMCӵ������崯,+�Ͱ�:��Y��^�ր�N�3O���y�,3O�_]L.�W��_�r[]H���E��������D���Q���^����=Ϸ�27����V#ol+���ҭ.�a�$ٷ_������'�+�:ʘ�a��U��_uJ��l?�f�O�H"nm�X7r�(�WH�K�˼B*]ǖ�8]1垣��2��M�Kj*�o��R�Ϥ�u�
��q�?a_מ���i�|9ў����Hq�$�}[$=L��2���uق95��	Zw�4����?o�yK�v�|�ݓa$�|l�_����Z�jy�?�_�.E_@k��U�Kh-Z�U���R��_�����l�B�s$��_���Ԓ�R=
]�ՇH�J�U)�*%V�Ī�X��RbUJ�J�Ui�\������šgB��Pu�6�6�1�����9-�㡓���W�oB߅.(�<��2�@��nS�j��ƨ	j�����\�����D��'X'g���U'}�F�U�^�~uPQ'�iuF�Sߪ�Տ�%��-x!b3�0G�w�c͉�Vəe����c�"�I�i�U+��*���dn7�0���a��j��q�k)�?X��X�֭� �ȹݺ�i�f�X9��`��Ul-f|X�v���}�\��e�h9�J^��SrzZ���*�,�
%�9��i��C�uՀ�Aע�������t#�*ڈ��nB7�M�t+�ݎ�@w��������^�-�}݇���G�E���C�a���=�E����я��'h+�)z=��F?C����v����V�Z]��0�ޖrŒ�>���>�����}����}��O\��\�+Pʀ_��D�^P6|�FP#�����S6|ʆO��)R�������<t6����Q�ѻ�1�=�Xt:^�H<������݂��%��]�}��>�xv~vָ�G�gg�򟊋��~U<��Is򋳳��.�3w��׷���W���
endstream
endobj
11 0 obj
<<
/BaseFont /CIDFont+F1
/DescendantFonts [ <<
/BaseFont /CIDFont+F1
/CIDSystemInfo <<
/Ordering 4 0 R
/Registry 5 0 R
/Supplement 0
>>
/CIDToGIDMap /Identity
/FontDescriptor <<
/Ascent 1000
/CapHeight 727
/Descent -206
/Flags 6
/FontBBox 6 0 R
/FontFile2 8 0 R
/FontName /CIDFont+F1
/ItalicAngle 0
/StemV 7 0 R
/Type /FontDescriptor
>>
/Subtype /CIDFontType2
/Type /Font
/W 9 0 R
>> ]
/Encoding /Identity-H
/Subtype /Type0
/ToUnicode 10 0 R
/Type /Font
>>
endobj
12 0 obj
<<
/Filter /FlateDecode
/Length 6721
>>
stream
x��O��Jv���)jm��+����{�/������0cL�����w�2�8G:��O@/ރ�WY�yu�
�h.�ؤ�^�K��?>�Mm���?�/��Ү������^�8_�6�8�vå����o�K3�G0����/ݜ�.&3����^���Ԃc�h���/���������k�~�����������C�A�ܛѾ~������f��-�b�B�F��~y�4��4}�:����M�6��m��m�O-kᷳV(O��~�Y�����ہ�1���������_~�~v������s���_�_��/�/�м�_
��B���/�cm�O�i�����7.E�<��	;\����J�pY�;&ɮ�/���8,�w4Om���]%c\�z�J�/K�L�����e�Ӷ���99&uMCv��:���i���Oݥ�CǍ(�F<��.s�;�	4ܻșà��|�H�0 �!��iw�}��XB(�0��B�|��_��k&�a:\6o��u�6���66?i�I���Mg��ӥ�8�������B9�`��|%F觷�HM^?��ݺJgМ�����'m{4}����8h����|��ff��4@�h/Ń��@�;���HNm�9�yYi�:�o��3o#g����"����O�vp}�>��r�vp�LWDj\�.>���O������4tM}|���o�9�߶�i�(�J����m';��K���o�r��W�pE�f��1�z{�(�f�4jЄڿUo������~�x��eM��z0��9L��q����^^�վ�}P)��-�m�gǤ+4��,��>n���)�� �{�F��|҈�a�Юg��`���f<� R1�r��̓yԬ\�G�͚7PT�m���m����Q�����I�Nb(�kNG1�.���%Q3�P�C@9����R.N~J-���0X�n������2���m,�66?i�ɸ���Hc(��C��"`��D*�R1��(�&�t�aZ�E��o^ټ��As�6���66?i�I�����bД�#M1S���A�CМ>c0���xr�\��;8�D����(�V��8�ʣ̮����x���l�e�,�ڶ��_g/t�87��I]�Y��d�k����d������)�6Y��I]�Y��d�8��҄,�̾T�W����.��T��G+�۾��d�����M�i\gf�<�K<�7�l����}@o�)Y�y})u���xyR�xVo*ٜgw��r+M���K�{�'4V��%�ӛR6Ӷ\�K�D3�R��p�##/O���M%{���JS�D��R�^�A��'u�g���M�a��#HY�y})uo�&�<�K<�7�l~8�/O�Z�S�D��R�^qZ�˓�ĳzS�&Zhj�R�h^_J�+>�5�����fT9BC�A���K�{}�y]�c�i]�9�)e��j�R�h^_J����*9��%�՛J6���Ҥ�&�ϝ�%�חR7�J��u�g���M����#HY�y})uoj��Z�xVo*�L�5r)K4�/���9\��:f��%�՛J6��\#G��D��R�&^��/{yR�xVo*�����z'M���K��xm_%GкĳzS�&Z�]�Ğ��N���K��x}��C���N���M%�hCS#G��D��R�f^�ti��E7O���M!�hc�4y����)Y�y})uo���Z�xVo*�D��KH#��|�,Ѽ�����*9��%�՛J6�b�7�ٻ�I���K�{}���A���M)�h	]!G��D��R�&^�\�tRg�\��%�՛J6��%��gg>wJ�hf_*��+ozyR�xVo*�D�9��%�חR7�ƱJ��u�g���M�iX��3M���K��x�u�
9��%�՛J6�BW#G��D��R�&^l�5���y��%�՛J6�b�A����(s��	Ur�K<�7�l��s�A���K��x�T%GкĳzS�&Z?�X�+e�����M�a��#h]�Y��dm�j�R�h^_J�ěڥ@p�;�K<�7�l��M�A���K��y��sz�K<�7�Z�0�P#G��D��R�&^����.��T�ח�L5V�JY�Y}�u/W���#h]�Y��d��k�R�h^_J���*ky�.��T��6�5r)K4�/�n�M���Z�xVo*�L�5r)K4�/�����Z�xVo*�D��+y�,Ѽ�����*9��%�՛J6��P#G��D��R�^_b�� �AM�X��I�O�t�9G��D��R�&^�� �AM�X��I�Ob.����,Ѽ������Z�x^oF�#�:A��+�;���J5A⃚ �Nœ�+��i��#HY�y})u�RM���&H�S�$�'�NE��+��J�N�z'�RM���&H�S�$�'mS�$��e�՝�b��(<f�٧Q�
mS�4��e�٣j��M.����(�������]��<]#�£'��ð<�K}�<nO�s�Ge'��M3����%�3�����P�t�aZ�6���v!6So��\2�y�*�^پ�~>rU�iy�p�C��W�,���K����I���+�ɇ�l4_��y+M��N^cڝ��T['ڝ�2�eڝ<�DN��#�B����q�
Jpov�uQ�bo��co��}�qS�ڝs2��Pp��PF�xd��JYz���+�;��Ƀ
�x����KC����>�;y�B���䕒e�C��W��1�Nm�x�G;�ԩ�;#S�܇�z�ю�0�T�s��_�s�2ehwG�����+����v#jk��N^)wEڭ�R�ڝ�R�yhw�J�&���[�����+u�8^����y`  ��0�%ۀ���	�N��1��y��:g�����vgp�BI�C��Wj1�N^�d&Bv#���ņv+�ܡ�Gv'���aڝ�R��yhw�f]��<�[y[����s{5}�뗔��sF;v¨S�sF̱s���
�pp��Ӽ��`ڝ�R��yhw�Rʦ2�;y��	_l`w���>�;ym[�B��v'�T�`ڭ�(3�;y�R��?�9O�6t��ؔ(t�h�Nu*vΈ9v��ꜧr�88���R
�yhw��Ց�v'���`ڝ�R��/6�[ye�t�}h�򢼹��ȃ��#��W*0�N^y5�����5mY6t�s�:g�c'�:;g�;��uιԀJ������?������v'���<�;y�u�����Eys%��W^�fڝ��5��n�����#��W�E�xA�G;���@ :��m���sF;v¨S�sF̱s��u��n5ڝ�Q^vfڝ���1�������v+/ʥQh���K�������X��v'��X�<�;ye�y��ȃ�/)^�ӥ�'�sT��˩d�9��:稧;ܝ3`���_�s��I)8����c�u���%��n�E�����+/%��v+����Xi�q,;�3�NރuǱҺ��r��D��䕷�8^����9�j�by�j,���t �aT��=#��=���g|y���m�U<��^�^~�����V�4�x�J,ou�uG�ļ�8�����F<`%��|�꼴�#%���;���eȈӫ������Y�� N� �>�D�~&j��G���NP!N�[YS.��L�:� �[�ࢢf9i������a}A�����߆�E�ZױCM¿�����'�/}nC�M:|_�~h(�?����}����m;��c�G�vN?;�.;t������[�Q#H����ؼEh�B��ww�_����[;��1����<
��hl�~�Ǚ�����žU;?��e��8���I�츅m�e���[�#m�9���c�︁��~x�_P��;�_��;O}8:�q���yN��u{#-��V?��^�����W��ʡ�׶4�J�e�*�wmϺ����q�'��ke�|M�����V1��9�C�"hv\ ʽ��e�m�槐���Yʩ���j�Q�_0s_���������׏5�~R��{�y����ʦy�2W��&������\���JV������)wïb���t{̙��w�@�z��$8x�1ޖf��1��� o�l�G=N��c� s� ����2�M���Ӵ��-�����ǔC��4�,f�i0�t�`L�4S:i0�D�)�4S"ƔN�)�cJ'ƔH�1��cJ����J+cJ��1���c����b�
�M���ќ/���"h�7��:����/KO7������3��j�1w��R=+?Ŏ��x[	j9�Ј�n��S#���'��-q�v�;����S3�o�@9������y�b8M���>���|䳷�CN!4Lǀ���3���F�U���'m;	�tc[tv�θ��LW�pE�f��1�{�(��+1B?�EGj�����3[kМ�����'m;)��l��0h��[�IǠ3F�T�|���-����ހ��#� +C{��~�F�d��΀;oEVi����$�`@�7�-���+f
�"R3�
�p��o~p�N��|od)�������Kր;mEVi����$�b�y	�4���㣀+f
�"R3�
�p�=h�O�c5h��C���
�l�(��+I�~} Ls��Ls����aP������t�Y��b�����3�>��M��+���욪ӏ�V�����:��4�~t�`�i0����#�`��I��G�����ӏH��G'��ӏNL?"���2�H�2�x����c.�0���Z<�/����{��\o�1�=/�i�����|��M�4�ѕ����Tl>.�K4槳ɱ�I7jD1�4�d6hh׳La0���xG3�o�H9��q9�yrH�8O�4[@��r{dsY�l��Q�����I�Nb(�0��e���1T�CE�f�,���cH��M,}W���"u��i�0X�ml~Ҷ���Խ��KkE[�!0c��H�B�!����i�����0:�H����cМ�������O�v4s)~�AS�G(h���������t�9���)��ءח���z+0J�h���L�zZcXW|�|K1�|Kޛ뾀�Dȼ�I]�sV M����t�1���i���y�ײ��Y�ڧ[�pvw�b�N� �L'�[��-NL� �[�4�nAL�8i0݂4�nq�`�i0���t�`��J+�-D+�-N$��MdWg��No������8����xyR�xVo*Y�c�J��wr�~+�}�o�r�<�K<�7�,��	Y��}�t�����{�u~�v��ț�����d����Խ�Ĺ�Ui�I]�Y��di�O+Mo������8�e���[�wj+��Yg��No������8�e_i�������ڿߊCo�^��%�ٗJ�68��l�߫}��8�f���Ҕ,Ѽ���W\��I]�Y��di�X+M���K�K�zyR�xVo*Y��JS�D��R�R�+/O���M%K��ZiJ�h^_J]��̋2G �כQ�����d����ԥ�~�<�K<�7�,�.l�)Y�y})ui/c/O���M%K;'[iJ�h^_J]ڧ�˓�ĳzS��v���#HY�y})u�V��'u�g����M����r0�}e� [D{yR�xVo*Yڐ�JS�D��R�޶���˓�ĳzS��f�N��%�՗Z�����.��T������d����ԥm˽<�K<�7��m��
9��%�חR�
m�yJ�x^o
Y���JS�D��R��ӧ*9��%�՛J��g�Ҕ,Ѽ������k�Z�xVo*Y�{�JS�D��R��N�V��%�ӛR���~�A���K�K��{yR�xVo*�L�μ^��%�ٗJ�v���.��T��-�+�R�h^_J���*9��%�՛J6Ѧaݷ�JS�D��R�&^~e�B��u�g���M�����,Ѽ�����mK +O���M%�i�F� e�f�e�9�܄*9��%�ӛR6�ڹF� e����ԥ-��<�K<�7�l��M��+y�,Ѽ����7Ur�K<�7�l��]�A���K��xS�m"d�I]�Y��dmnj�R�h^_J�̋U��k]�y��*�9�9��%�חR7��F��u�g������f���W���K�K��zyR�xVo*�D��9��%�חR7����Z^�K<�7�l�m�A���K��xcSe-��%�՛J6�b�A����(s�0�*9��%�՛J6���J^)K4�/�nⅱJ��u�g���M�8���,Ѽ���������u*�D]�$�Kw�s)K4�/�n�U�	��u*�D]�$���A���K��y�J��u���fT9B�S$� �R�����I�T$>�	�T<���I��9��%�חR7�*��j��:O��x�T��"H�T�$>�w+��j��:O��x�6uJ�h]�Y��@x!�*��a&�}U��6uJ�h]�=���I��B��8��R��^�*]����5B�.<�����a���+��`'{����a>�ݛ| e�}��w�����">Tn�ã#�n������3�s��oGf��]��';�7Ka�\��������Owm���T�Yjڏ��n�2ʻ_�/�����e���o��^��b,ϼ+(�o�b����nG.n0o�5Ʒ�ű��b.���_�����-���g��Z�+Z��w�t��w&{y�&�K��sS�=�=�9�Z��q��ݶ������~�ȗÁm��{j��Pl��g�i���fwEӹ����M�:�]#ڷ�z�b�/�B�7�۷b9�z1�5�ڟ�ݦ��}S�r������r�O��.�w�m�͟ί!�x�,_�8���>����U��o	��b8�I
endstream
endobj
13 0 obj
<<
/Font <<
/F1 11 0 R
>>
>>
endobj
3 0 obj
<<
/Contents [ 12 0 R ]
/CropBox [ 0.0 0.0 792.0 612.0 ]
/MediaBox [ 0.0 0.0 792.0 612.0 ]
/Parent 2 0 R
/Resources 13 0 R
/Rotate 0
/Type /Page
>>
endobj
10 0 obj
<<
/Length 969
>>
stream
/CIDInit /ProcSet findresource begin 12 dict begin begincmap /CIDSystemInfo << /Registry (Adobe) /Ordering (UCS) /Supplement 0 >> def /CMapName /Adobe-Identity-UCS def /CMapType 2 def 1 begincodespacerange <0000> <FFFF> endcodespacerange 46 beginbfchar <0003> <0020> <0012> <002F> <0013> <0030> <0014> <0031> <0015> <0032> <0016> <0033> <0017> <0034> <0018> <0035> <0019> <0036> <001A> <0037> <001B> <0038> <001C> <0039> <001D> <003A> <0024> <0041> <0027> <0044> <0028> <0045> <0030> <004D> <0031> <004E> <0033> <0050> <0035> <0052> <0036> <0053> <0037> <0054> <003B> <0058> <0042> <005F> <0044> <0061> <0045> <0062> <0046> <0063> <0047> <0064> <0048> <0065> <004A> <0067> <004B> <0068> <004C> <0069> <004E> <006B> <004F> <006C> <0050> <006D> <0051> <006E> <0052> <006F> <0055> <0072> <0056> <0073> <0057> <0074> <0058> <0075> <0059> <0076> <005A> <0077> <005C> <0079> <005E> <007B> <0060> <007D> endbfchar endcmap CMapName currentdict /CMap defineresource pop end end 
endstream
endobj
9 0 obj
[ 3 3 312 18 18 382 19 19 545 20 20 545 21 21 545 22 22 545 23 23 545 24 24 545 25 25 545 26 26 545 27 27 545 28 28 545 29 29 353 36 36 599 39 39 678 40 40 561 48 48 770 49 49 667 51 51 551 53 53 620 54 54 557 55 55 583 59 59 580 66 66 545 68 68 524 69 69 552 70 70 461 71 71 552 72 72 526 74 74 552 75 75 557 76 76 228 78 78 498 79 79 228 80 80 839 81 81 557 82 82 542 85 85 360 86 86 446 87 87 334 88 88 557 89 89 498 90 90 742 92 92 498 94 94 480 96 96 480 ]
endobj
6 0 obj
[ -839 -206 839 1000 ]
endobj
7 0 obj
839
endobj
2 0 obj
<<
/Count 1
/Kids [ 3 0 R ]
/Type /Pages
>>
endobj
1 0 obj
<<
/Pages 2 0 R
/Type /Catalog
>>
endobj
14 0 obj
<<
/Author (martinda3)
/CreationDate (D:20191111083753-05'00')
/ModDate (D:20191111083753-05'00')
/Producer (Microsoft: Print To PDF)
/Title (ModelSim: instruction_mem_tb(behavioral))
>>
endobj
xref
0 15
0000000000 65535 f
0000076258 00000 n
0000076199 00000 n
0000074481 00000 n
0000000009 00000 n
0000000035 00000 n
0000076142 00000 n
0000076180 00000 n
0000000058 00000 n
0000075665 00000 n
0000074644 00000 n
0000067168 00000 n
0000067641 00000 n
0000074436 00000 n
0000076307 00000 n
trailer
<<
/Info 14 0 R
/Root 1 0 R
/Size 15
>>
startxref
76511
%%EOF
